//==========================================================
//      RTL Generated File
//      Author: Ashish Tondwalkar
//--------------------------------------------------
//      Description: Systolic Array of MAC Units
//--------------------------------------------------
//      Datawidth = 16
//      Dimension = 32
//==========================================================

module ast_systolic_array_v (
    a_in,
    b_in,
    mult_en,
    acc_en,
    load_en,
    clk,
    reset,
    d_out,
    );

    localparam DATAWIDTH = 15;
    localparam SIZE = 31;

    input clk, reset, mult_en, acc_en, load_en;
    input [DATAWIDTH:0] a_in [SIZE:0]; //data input from row fifo set
    input [DATAWIDTH:0] b_in [SIZE:0]; //data input from col fifo set
    output reg  [SIZE:0][SIZE:0][DATAWIDTH:0] d_out;

    wire [SIZE+1:0][SIZE+1:0][DATAWIDTH:0] a; //internal array row connections
    wire [SIZE+1:0][SIZE+1:0][DATAWIDTH:0] b; //internal array col connections


    //row bounday
    assign a[0][0] = a_in[0];
    assign a[1][0] = a_in[1];
    assign a[2][0] = a_in[2];
    assign a[3][0] = a_in[3];
    assign a[4][0] = a_in[4];
    assign a[5][0] = a_in[5];
    assign a[6][0] = a_in[6];
    assign a[7][0] = a_in[7];
    assign a[8][0] = a_in[8];
    assign a[9][0] = a_in[9];
    assign a[10][0] = a_in[10];
    assign a[11][0] = a_in[11];
    assign a[12][0] = a_in[12];
    assign a[13][0] = a_in[13];
    assign a[14][0] = a_in[14];
    assign a[15][0] = a_in[15];
    assign a[16][0] = a_in[16];
    assign a[17][0] = a_in[17];
    assign a[18][0] = a_in[18];
    assign a[19][0] = a_in[19];
    assign a[20][0] = a_in[20];
    assign a[21][0] = a_in[21];
    assign a[22][0] = a_in[22];
    assign a[23][0] = a_in[23];
    assign a[24][0] = a_in[24];
    assign a[25][0] = a_in[25];
    assign a[26][0] = a_in[26];
    assign a[27][0] = a_in[27];
    assign a[28][0] = a_in[28];
    assign a[29][0] = a_in[29];
    assign a[30][0] = a_in[30];
    assign a[31][0] = a_in[31];

    //col bounday
    assign b[0][0] = b_in[0];
    assign b[0][1] = b_in[1];
    assign b[0][2] = b_in[2];
    assign b[0][3] = b_in[3];
    assign b[0][4] = b_in[4];
    assign b[0][5] = b_in[5];
    assign b[0][6] = b_in[6];
    assign b[0][7] = b_in[7];
    assign b[0][8] = b_in[8];
    assign b[0][9] = b_in[9];
    assign b[0][10] = b_in[10];
    assign b[0][11] = b_in[11];
    assign b[0][12] = b_in[12];
    assign b[0][13] = b_in[13];
    assign b[0][14] = b_in[14];
    assign b[0][15] = b_in[15];
    assign b[0][16] = b_in[16];
    assign b[0][17] = b_in[17];
    assign b[0][18] = b_in[18];
    assign b[0][19] = b_in[19];
    assign b[0][20] = b_in[20];
    assign b[0][21] = b_in[21];
    assign b[0][22] = b_in[22];
    assign b[0][23] = b_in[23];
    assign b[0][24] = b_in[24];
    assign b[0][25] = b_in[25];
    assign b[0][26] = b_in[26];
    assign b[0][27] = b_in[27];
    assign b[0][28] = b_in[28];
    assign b[0][29] = b_in[29];
    assign b[0][30] = b_in[30];
    assign b[0][31] = b_in[31];

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][0]), 
        .b_in(b[0][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][1]), 
        .b_out(b[1][0]),
        .acc_out(d_out[0][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][1]), 
        .b_in(b[0][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][2]), 
        .b_out(b[1][1]),
        .acc_out(d_out[0][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][2]), 
        .b_in(b[0][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][3]), 
        .b_out(b[1][2]),
        .acc_out(d_out[0][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][3]), 
        .b_in(b[0][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][4]), 
        .b_out(b[1][3]),
        .acc_out(d_out[0][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][4]), 
        .b_in(b[0][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][5]), 
        .b_out(b[1][4]),
        .acc_out(d_out[0][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][5]), 
        .b_in(b[0][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][6]), 
        .b_out(b[1][5]),
        .acc_out(d_out[0][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][6]), 
        .b_in(b[0][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][7]), 
        .b_out(b[1][6]),
        .acc_out(d_out[0][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][7]), 
        .b_in(b[0][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][8]), 
        .b_out(b[1][7]),
        .acc_out(d_out[0][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][8]), 
        .b_in(b[0][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][9]), 
        .b_out(b[1][8]),
        .acc_out(d_out[0][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][9]), 
        .b_in(b[0][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][10]), 
        .b_out(b[1][9]),
        .acc_out(d_out[0][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][10]), 
        .b_in(b[0][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][11]), 
        .b_out(b[1][10]),
        .acc_out(d_out[0][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][11]), 
        .b_in(b[0][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][12]), 
        .b_out(b[1][11]),
        .acc_out(d_out[0][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][12]), 
        .b_in(b[0][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][13]), 
        .b_out(b[1][12]),
        .acc_out(d_out[0][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][13]), 
        .b_in(b[0][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][14]), 
        .b_out(b[1][13]),
        .acc_out(d_out[0][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][14]), 
        .b_in(b[0][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][15]), 
        .b_out(b[1][14]),
        .acc_out(d_out[0][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][15]), 
        .b_in(b[0][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][16]), 
        .b_out(b[1][15]),
        .acc_out(d_out[0][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][16]), 
        .b_in(b[0][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][17]), 
        .b_out(b[1][16]),
        .acc_out(d_out[0][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][17]), 
        .b_in(b[0][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][18]), 
        .b_out(b[1][17]),
        .acc_out(d_out[0][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][18]), 
        .b_in(b[0][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][19]), 
        .b_out(b[1][18]),
        .acc_out(d_out[0][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][19]), 
        .b_in(b[0][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][20]), 
        .b_out(b[1][19]),
        .acc_out(d_out[0][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][20]), 
        .b_in(b[0][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][21]), 
        .b_out(b[1][20]),
        .acc_out(d_out[0][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][21]), 
        .b_in(b[0][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][22]), 
        .b_out(b[1][21]),
        .acc_out(d_out[0][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][22]), 
        .b_in(b[0][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][23]), 
        .b_out(b[1][22]),
        .acc_out(d_out[0][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][23]), 
        .b_in(b[0][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][24]), 
        .b_out(b[1][23]),
        .acc_out(d_out[0][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][24]), 
        .b_in(b[0][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][25]), 
        .b_out(b[1][24]),
        .acc_out(d_out[0][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][25]), 
        .b_in(b[0][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][26]), 
        .b_out(b[1][25]),
        .acc_out(d_out[0][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][26]), 
        .b_in(b[0][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][27]), 
        .b_out(b[1][26]),
        .acc_out(d_out[0][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][27]), 
        .b_in(b[0][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][28]), 
        .b_out(b[1][27]),
        .acc_out(d_out[0][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][28]), 
        .b_in(b[0][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][29]), 
        .b_out(b[1][28]),
        .acc_out(d_out[0][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][29]), 
        .b_in(b[0][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][30]), 
        .b_out(b[1][29]),
        .acc_out(d_out[0][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][30]), 
        .b_in(b[0][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][31]), 
        .b_out(b[1][30]),
        .acc_out(d_out[0][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[0][31]), 
        .b_in(b[0][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[0][32]), 
        .b_out(b[1][31]),
        .acc_out(d_out[0][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][0]), 
        .b_in(b[1][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][1]), 
        .b_out(b[2][0]),
        .acc_out(d_out[1][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][1]), 
        .b_in(b[1][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][2]), 
        .b_out(b[2][1]),
        .acc_out(d_out[1][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][2]), 
        .b_in(b[1][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][3]), 
        .b_out(b[2][2]),
        .acc_out(d_out[1][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][3]), 
        .b_in(b[1][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][4]), 
        .b_out(b[2][3]),
        .acc_out(d_out[1][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][4]), 
        .b_in(b[1][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][5]), 
        .b_out(b[2][4]),
        .acc_out(d_out[1][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][5]), 
        .b_in(b[1][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][6]), 
        .b_out(b[2][5]),
        .acc_out(d_out[1][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][6]), 
        .b_in(b[1][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][7]), 
        .b_out(b[2][6]),
        .acc_out(d_out[1][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][7]), 
        .b_in(b[1][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][8]), 
        .b_out(b[2][7]),
        .acc_out(d_out[1][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][8]), 
        .b_in(b[1][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][9]), 
        .b_out(b[2][8]),
        .acc_out(d_out[1][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][9]), 
        .b_in(b[1][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][10]), 
        .b_out(b[2][9]),
        .acc_out(d_out[1][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][10]), 
        .b_in(b[1][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][11]), 
        .b_out(b[2][10]),
        .acc_out(d_out[1][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][11]), 
        .b_in(b[1][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][12]), 
        .b_out(b[2][11]),
        .acc_out(d_out[1][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][12]), 
        .b_in(b[1][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][13]), 
        .b_out(b[2][12]),
        .acc_out(d_out[1][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][13]), 
        .b_in(b[1][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][14]), 
        .b_out(b[2][13]),
        .acc_out(d_out[1][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][14]), 
        .b_in(b[1][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][15]), 
        .b_out(b[2][14]),
        .acc_out(d_out[1][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][15]), 
        .b_in(b[1][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][16]), 
        .b_out(b[2][15]),
        .acc_out(d_out[1][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][16]), 
        .b_in(b[1][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][17]), 
        .b_out(b[2][16]),
        .acc_out(d_out[1][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][17]), 
        .b_in(b[1][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][18]), 
        .b_out(b[2][17]),
        .acc_out(d_out[1][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][18]), 
        .b_in(b[1][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][19]), 
        .b_out(b[2][18]),
        .acc_out(d_out[1][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][19]), 
        .b_in(b[1][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][20]), 
        .b_out(b[2][19]),
        .acc_out(d_out[1][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][20]), 
        .b_in(b[1][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][21]), 
        .b_out(b[2][20]),
        .acc_out(d_out[1][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][21]), 
        .b_in(b[1][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][22]), 
        .b_out(b[2][21]),
        .acc_out(d_out[1][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][22]), 
        .b_in(b[1][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][23]), 
        .b_out(b[2][22]),
        .acc_out(d_out[1][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][23]), 
        .b_in(b[1][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][24]), 
        .b_out(b[2][23]),
        .acc_out(d_out[1][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][24]), 
        .b_in(b[1][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][25]), 
        .b_out(b[2][24]),
        .acc_out(d_out[1][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][25]), 
        .b_in(b[1][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][26]), 
        .b_out(b[2][25]),
        .acc_out(d_out[1][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][26]), 
        .b_in(b[1][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][27]), 
        .b_out(b[2][26]),
        .acc_out(d_out[1][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][27]), 
        .b_in(b[1][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][28]), 
        .b_out(b[2][27]),
        .acc_out(d_out[1][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][28]), 
        .b_in(b[1][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][29]), 
        .b_out(b[2][28]),
        .acc_out(d_out[1][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][29]), 
        .b_in(b[1][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][30]), 
        .b_out(b[2][29]),
        .acc_out(d_out[1][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][30]), 
        .b_in(b[1][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][31]), 
        .b_out(b[2][30]),
        .acc_out(d_out[1][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[1][31]), 
        .b_in(b[1][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[1][32]), 
        .b_out(b[2][31]),
        .acc_out(d_out[1][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][0]), 
        .b_in(b[2][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][1]), 
        .b_out(b[3][0]),
        .acc_out(d_out[2][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][1]), 
        .b_in(b[2][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][2]), 
        .b_out(b[3][1]),
        .acc_out(d_out[2][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][2]), 
        .b_in(b[2][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][3]), 
        .b_out(b[3][2]),
        .acc_out(d_out[2][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][3]), 
        .b_in(b[2][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][4]), 
        .b_out(b[3][3]),
        .acc_out(d_out[2][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][4]), 
        .b_in(b[2][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][5]), 
        .b_out(b[3][4]),
        .acc_out(d_out[2][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][5]), 
        .b_in(b[2][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][6]), 
        .b_out(b[3][5]),
        .acc_out(d_out[2][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][6]), 
        .b_in(b[2][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][7]), 
        .b_out(b[3][6]),
        .acc_out(d_out[2][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][7]), 
        .b_in(b[2][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][8]), 
        .b_out(b[3][7]),
        .acc_out(d_out[2][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][8]), 
        .b_in(b[2][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][9]), 
        .b_out(b[3][8]),
        .acc_out(d_out[2][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][9]), 
        .b_in(b[2][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][10]), 
        .b_out(b[3][9]),
        .acc_out(d_out[2][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][10]), 
        .b_in(b[2][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][11]), 
        .b_out(b[3][10]),
        .acc_out(d_out[2][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][11]), 
        .b_in(b[2][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][12]), 
        .b_out(b[3][11]),
        .acc_out(d_out[2][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][12]), 
        .b_in(b[2][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][13]), 
        .b_out(b[3][12]),
        .acc_out(d_out[2][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][13]), 
        .b_in(b[2][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][14]), 
        .b_out(b[3][13]),
        .acc_out(d_out[2][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][14]), 
        .b_in(b[2][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][15]), 
        .b_out(b[3][14]),
        .acc_out(d_out[2][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][15]), 
        .b_in(b[2][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][16]), 
        .b_out(b[3][15]),
        .acc_out(d_out[2][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][16]), 
        .b_in(b[2][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][17]), 
        .b_out(b[3][16]),
        .acc_out(d_out[2][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][17]), 
        .b_in(b[2][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][18]), 
        .b_out(b[3][17]),
        .acc_out(d_out[2][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][18]), 
        .b_in(b[2][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][19]), 
        .b_out(b[3][18]),
        .acc_out(d_out[2][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][19]), 
        .b_in(b[2][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][20]), 
        .b_out(b[3][19]),
        .acc_out(d_out[2][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][20]), 
        .b_in(b[2][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][21]), 
        .b_out(b[3][20]),
        .acc_out(d_out[2][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][21]), 
        .b_in(b[2][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][22]), 
        .b_out(b[3][21]),
        .acc_out(d_out[2][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][22]), 
        .b_in(b[2][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][23]), 
        .b_out(b[3][22]),
        .acc_out(d_out[2][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][23]), 
        .b_in(b[2][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][24]), 
        .b_out(b[3][23]),
        .acc_out(d_out[2][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][24]), 
        .b_in(b[2][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][25]), 
        .b_out(b[3][24]),
        .acc_out(d_out[2][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][25]), 
        .b_in(b[2][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][26]), 
        .b_out(b[3][25]),
        .acc_out(d_out[2][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][26]), 
        .b_in(b[2][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][27]), 
        .b_out(b[3][26]),
        .acc_out(d_out[2][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][27]), 
        .b_in(b[2][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][28]), 
        .b_out(b[3][27]),
        .acc_out(d_out[2][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][28]), 
        .b_in(b[2][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][29]), 
        .b_out(b[3][28]),
        .acc_out(d_out[2][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][29]), 
        .b_in(b[2][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][30]), 
        .b_out(b[3][29]),
        .acc_out(d_out[2][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][30]), 
        .b_in(b[2][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][31]), 
        .b_out(b[3][30]),
        .acc_out(d_out[2][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[2][31]), 
        .b_in(b[2][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[2][32]), 
        .b_out(b[3][31]),
        .acc_out(d_out[2][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][0]), 
        .b_in(b[3][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][1]), 
        .b_out(b[4][0]),
        .acc_out(d_out[3][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][1]), 
        .b_in(b[3][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][2]), 
        .b_out(b[4][1]),
        .acc_out(d_out[3][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][2]), 
        .b_in(b[3][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][3]), 
        .b_out(b[4][2]),
        .acc_out(d_out[3][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][3]), 
        .b_in(b[3][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][4]), 
        .b_out(b[4][3]),
        .acc_out(d_out[3][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][4]), 
        .b_in(b[3][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][5]), 
        .b_out(b[4][4]),
        .acc_out(d_out[3][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][5]), 
        .b_in(b[3][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][6]), 
        .b_out(b[4][5]),
        .acc_out(d_out[3][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][6]), 
        .b_in(b[3][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][7]), 
        .b_out(b[4][6]),
        .acc_out(d_out[3][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][7]), 
        .b_in(b[3][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][8]), 
        .b_out(b[4][7]),
        .acc_out(d_out[3][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][8]), 
        .b_in(b[3][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][9]), 
        .b_out(b[4][8]),
        .acc_out(d_out[3][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][9]), 
        .b_in(b[3][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][10]), 
        .b_out(b[4][9]),
        .acc_out(d_out[3][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][10]), 
        .b_in(b[3][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][11]), 
        .b_out(b[4][10]),
        .acc_out(d_out[3][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][11]), 
        .b_in(b[3][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][12]), 
        .b_out(b[4][11]),
        .acc_out(d_out[3][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][12]), 
        .b_in(b[3][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][13]), 
        .b_out(b[4][12]),
        .acc_out(d_out[3][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][13]), 
        .b_in(b[3][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][14]), 
        .b_out(b[4][13]),
        .acc_out(d_out[3][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][14]), 
        .b_in(b[3][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][15]), 
        .b_out(b[4][14]),
        .acc_out(d_out[3][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][15]), 
        .b_in(b[3][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][16]), 
        .b_out(b[4][15]),
        .acc_out(d_out[3][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][16]), 
        .b_in(b[3][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][17]), 
        .b_out(b[4][16]),
        .acc_out(d_out[3][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][17]), 
        .b_in(b[3][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][18]), 
        .b_out(b[4][17]),
        .acc_out(d_out[3][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][18]), 
        .b_in(b[3][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][19]), 
        .b_out(b[4][18]),
        .acc_out(d_out[3][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][19]), 
        .b_in(b[3][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][20]), 
        .b_out(b[4][19]),
        .acc_out(d_out[3][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][20]), 
        .b_in(b[3][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][21]), 
        .b_out(b[4][20]),
        .acc_out(d_out[3][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][21]), 
        .b_in(b[3][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][22]), 
        .b_out(b[4][21]),
        .acc_out(d_out[3][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][22]), 
        .b_in(b[3][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][23]), 
        .b_out(b[4][22]),
        .acc_out(d_out[3][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][23]), 
        .b_in(b[3][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][24]), 
        .b_out(b[4][23]),
        .acc_out(d_out[3][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][24]), 
        .b_in(b[3][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][25]), 
        .b_out(b[4][24]),
        .acc_out(d_out[3][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][25]), 
        .b_in(b[3][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][26]), 
        .b_out(b[4][25]),
        .acc_out(d_out[3][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][26]), 
        .b_in(b[3][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][27]), 
        .b_out(b[4][26]),
        .acc_out(d_out[3][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][27]), 
        .b_in(b[3][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][28]), 
        .b_out(b[4][27]),
        .acc_out(d_out[3][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][28]), 
        .b_in(b[3][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][29]), 
        .b_out(b[4][28]),
        .acc_out(d_out[3][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][29]), 
        .b_in(b[3][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][30]), 
        .b_out(b[4][29]),
        .acc_out(d_out[3][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][30]), 
        .b_in(b[3][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][31]), 
        .b_out(b[4][30]),
        .acc_out(d_out[3][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[3][31]), 
        .b_in(b[3][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[3][32]), 
        .b_out(b[4][31]),
        .acc_out(d_out[3][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][0]), 
        .b_in(b[4][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][1]), 
        .b_out(b[5][0]),
        .acc_out(d_out[4][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][1]), 
        .b_in(b[4][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][2]), 
        .b_out(b[5][1]),
        .acc_out(d_out[4][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][2]), 
        .b_in(b[4][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][3]), 
        .b_out(b[5][2]),
        .acc_out(d_out[4][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][3]), 
        .b_in(b[4][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][4]), 
        .b_out(b[5][3]),
        .acc_out(d_out[4][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][4]), 
        .b_in(b[4][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][5]), 
        .b_out(b[5][4]),
        .acc_out(d_out[4][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][5]), 
        .b_in(b[4][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][6]), 
        .b_out(b[5][5]),
        .acc_out(d_out[4][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][6]), 
        .b_in(b[4][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][7]), 
        .b_out(b[5][6]),
        .acc_out(d_out[4][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][7]), 
        .b_in(b[4][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][8]), 
        .b_out(b[5][7]),
        .acc_out(d_out[4][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][8]), 
        .b_in(b[4][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][9]), 
        .b_out(b[5][8]),
        .acc_out(d_out[4][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][9]), 
        .b_in(b[4][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][10]), 
        .b_out(b[5][9]),
        .acc_out(d_out[4][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][10]), 
        .b_in(b[4][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][11]), 
        .b_out(b[5][10]),
        .acc_out(d_out[4][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][11]), 
        .b_in(b[4][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][12]), 
        .b_out(b[5][11]),
        .acc_out(d_out[4][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][12]), 
        .b_in(b[4][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][13]), 
        .b_out(b[5][12]),
        .acc_out(d_out[4][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][13]), 
        .b_in(b[4][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][14]), 
        .b_out(b[5][13]),
        .acc_out(d_out[4][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][14]), 
        .b_in(b[4][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][15]), 
        .b_out(b[5][14]),
        .acc_out(d_out[4][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][15]), 
        .b_in(b[4][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][16]), 
        .b_out(b[5][15]),
        .acc_out(d_out[4][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][16]), 
        .b_in(b[4][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][17]), 
        .b_out(b[5][16]),
        .acc_out(d_out[4][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][17]), 
        .b_in(b[4][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][18]), 
        .b_out(b[5][17]),
        .acc_out(d_out[4][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][18]), 
        .b_in(b[4][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][19]), 
        .b_out(b[5][18]),
        .acc_out(d_out[4][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][19]), 
        .b_in(b[4][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][20]), 
        .b_out(b[5][19]),
        .acc_out(d_out[4][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][20]), 
        .b_in(b[4][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][21]), 
        .b_out(b[5][20]),
        .acc_out(d_out[4][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][21]), 
        .b_in(b[4][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][22]), 
        .b_out(b[5][21]),
        .acc_out(d_out[4][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][22]), 
        .b_in(b[4][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][23]), 
        .b_out(b[5][22]),
        .acc_out(d_out[4][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][23]), 
        .b_in(b[4][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][24]), 
        .b_out(b[5][23]),
        .acc_out(d_out[4][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][24]), 
        .b_in(b[4][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][25]), 
        .b_out(b[5][24]),
        .acc_out(d_out[4][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][25]), 
        .b_in(b[4][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][26]), 
        .b_out(b[5][25]),
        .acc_out(d_out[4][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][26]), 
        .b_in(b[4][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][27]), 
        .b_out(b[5][26]),
        .acc_out(d_out[4][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][27]), 
        .b_in(b[4][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][28]), 
        .b_out(b[5][27]),
        .acc_out(d_out[4][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][28]), 
        .b_in(b[4][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][29]), 
        .b_out(b[5][28]),
        .acc_out(d_out[4][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][29]), 
        .b_in(b[4][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][30]), 
        .b_out(b[5][29]),
        .acc_out(d_out[4][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][30]), 
        .b_in(b[4][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][31]), 
        .b_out(b[5][30]),
        .acc_out(d_out[4][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[4][31]), 
        .b_in(b[4][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[4][32]), 
        .b_out(b[5][31]),
        .acc_out(d_out[4][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][0]), 
        .b_in(b[5][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][1]), 
        .b_out(b[6][0]),
        .acc_out(d_out[5][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][1]), 
        .b_in(b[5][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][2]), 
        .b_out(b[6][1]),
        .acc_out(d_out[5][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][2]), 
        .b_in(b[5][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][3]), 
        .b_out(b[6][2]),
        .acc_out(d_out[5][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][3]), 
        .b_in(b[5][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][4]), 
        .b_out(b[6][3]),
        .acc_out(d_out[5][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][4]), 
        .b_in(b[5][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][5]), 
        .b_out(b[6][4]),
        .acc_out(d_out[5][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][5]), 
        .b_in(b[5][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][6]), 
        .b_out(b[6][5]),
        .acc_out(d_out[5][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][6]), 
        .b_in(b[5][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][7]), 
        .b_out(b[6][6]),
        .acc_out(d_out[5][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][7]), 
        .b_in(b[5][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][8]), 
        .b_out(b[6][7]),
        .acc_out(d_out[5][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][8]), 
        .b_in(b[5][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][9]), 
        .b_out(b[6][8]),
        .acc_out(d_out[5][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][9]), 
        .b_in(b[5][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][10]), 
        .b_out(b[6][9]),
        .acc_out(d_out[5][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][10]), 
        .b_in(b[5][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][11]), 
        .b_out(b[6][10]),
        .acc_out(d_out[5][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][11]), 
        .b_in(b[5][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][12]), 
        .b_out(b[6][11]),
        .acc_out(d_out[5][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][12]), 
        .b_in(b[5][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][13]), 
        .b_out(b[6][12]),
        .acc_out(d_out[5][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][13]), 
        .b_in(b[5][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][14]), 
        .b_out(b[6][13]),
        .acc_out(d_out[5][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][14]), 
        .b_in(b[5][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][15]), 
        .b_out(b[6][14]),
        .acc_out(d_out[5][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][15]), 
        .b_in(b[5][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][16]), 
        .b_out(b[6][15]),
        .acc_out(d_out[5][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][16]), 
        .b_in(b[5][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][17]), 
        .b_out(b[6][16]),
        .acc_out(d_out[5][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][17]), 
        .b_in(b[5][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][18]), 
        .b_out(b[6][17]),
        .acc_out(d_out[5][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][18]), 
        .b_in(b[5][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][19]), 
        .b_out(b[6][18]),
        .acc_out(d_out[5][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][19]), 
        .b_in(b[5][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][20]), 
        .b_out(b[6][19]),
        .acc_out(d_out[5][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][20]), 
        .b_in(b[5][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][21]), 
        .b_out(b[6][20]),
        .acc_out(d_out[5][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][21]), 
        .b_in(b[5][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][22]), 
        .b_out(b[6][21]),
        .acc_out(d_out[5][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][22]), 
        .b_in(b[5][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][23]), 
        .b_out(b[6][22]),
        .acc_out(d_out[5][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][23]), 
        .b_in(b[5][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][24]), 
        .b_out(b[6][23]),
        .acc_out(d_out[5][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][24]), 
        .b_in(b[5][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][25]), 
        .b_out(b[6][24]),
        .acc_out(d_out[5][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][25]), 
        .b_in(b[5][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][26]), 
        .b_out(b[6][25]),
        .acc_out(d_out[5][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][26]), 
        .b_in(b[5][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][27]), 
        .b_out(b[6][26]),
        .acc_out(d_out[5][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][27]), 
        .b_in(b[5][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][28]), 
        .b_out(b[6][27]),
        .acc_out(d_out[5][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][28]), 
        .b_in(b[5][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][29]), 
        .b_out(b[6][28]),
        .acc_out(d_out[5][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][29]), 
        .b_in(b[5][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][30]), 
        .b_out(b[6][29]),
        .acc_out(d_out[5][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][30]), 
        .b_in(b[5][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][31]), 
        .b_out(b[6][30]),
        .acc_out(d_out[5][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[5][31]), 
        .b_in(b[5][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[5][32]), 
        .b_out(b[6][31]),
        .acc_out(d_out[5][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][0]), 
        .b_in(b[6][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][1]), 
        .b_out(b[7][0]),
        .acc_out(d_out[6][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][1]), 
        .b_in(b[6][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][2]), 
        .b_out(b[7][1]),
        .acc_out(d_out[6][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][2]), 
        .b_in(b[6][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][3]), 
        .b_out(b[7][2]),
        .acc_out(d_out[6][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][3]), 
        .b_in(b[6][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][4]), 
        .b_out(b[7][3]),
        .acc_out(d_out[6][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][4]), 
        .b_in(b[6][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][5]), 
        .b_out(b[7][4]),
        .acc_out(d_out[6][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][5]), 
        .b_in(b[6][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][6]), 
        .b_out(b[7][5]),
        .acc_out(d_out[6][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][6]), 
        .b_in(b[6][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][7]), 
        .b_out(b[7][6]),
        .acc_out(d_out[6][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][7]), 
        .b_in(b[6][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][8]), 
        .b_out(b[7][7]),
        .acc_out(d_out[6][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][8]), 
        .b_in(b[6][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][9]), 
        .b_out(b[7][8]),
        .acc_out(d_out[6][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][9]), 
        .b_in(b[6][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][10]), 
        .b_out(b[7][9]),
        .acc_out(d_out[6][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][10]), 
        .b_in(b[6][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][11]), 
        .b_out(b[7][10]),
        .acc_out(d_out[6][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][11]), 
        .b_in(b[6][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][12]), 
        .b_out(b[7][11]),
        .acc_out(d_out[6][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][12]), 
        .b_in(b[6][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][13]), 
        .b_out(b[7][12]),
        .acc_out(d_out[6][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][13]), 
        .b_in(b[6][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][14]), 
        .b_out(b[7][13]),
        .acc_out(d_out[6][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][14]), 
        .b_in(b[6][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][15]), 
        .b_out(b[7][14]),
        .acc_out(d_out[6][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][15]), 
        .b_in(b[6][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][16]), 
        .b_out(b[7][15]),
        .acc_out(d_out[6][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][16]), 
        .b_in(b[6][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][17]), 
        .b_out(b[7][16]),
        .acc_out(d_out[6][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][17]), 
        .b_in(b[6][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][18]), 
        .b_out(b[7][17]),
        .acc_out(d_out[6][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][18]), 
        .b_in(b[6][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][19]), 
        .b_out(b[7][18]),
        .acc_out(d_out[6][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][19]), 
        .b_in(b[6][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][20]), 
        .b_out(b[7][19]),
        .acc_out(d_out[6][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][20]), 
        .b_in(b[6][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][21]), 
        .b_out(b[7][20]),
        .acc_out(d_out[6][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][21]), 
        .b_in(b[6][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][22]), 
        .b_out(b[7][21]),
        .acc_out(d_out[6][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][22]), 
        .b_in(b[6][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][23]), 
        .b_out(b[7][22]),
        .acc_out(d_out[6][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][23]), 
        .b_in(b[6][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][24]), 
        .b_out(b[7][23]),
        .acc_out(d_out[6][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][24]), 
        .b_in(b[6][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][25]), 
        .b_out(b[7][24]),
        .acc_out(d_out[6][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][25]), 
        .b_in(b[6][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][26]), 
        .b_out(b[7][25]),
        .acc_out(d_out[6][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][26]), 
        .b_in(b[6][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][27]), 
        .b_out(b[7][26]),
        .acc_out(d_out[6][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][27]), 
        .b_in(b[6][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][28]), 
        .b_out(b[7][27]),
        .acc_out(d_out[6][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][28]), 
        .b_in(b[6][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][29]), 
        .b_out(b[7][28]),
        .acc_out(d_out[6][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][29]), 
        .b_in(b[6][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][30]), 
        .b_out(b[7][29]),
        .acc_out(d_out[6][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][30]), 
        .b_in(b[6][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][31]), 
        .b_out(b[7][30]),
        .acc_out(d_out[6][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[6][31]), 
        .b_in(b[6][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[6][32]), 
        .b_out(b[7][31]),
        .acc_out(d_out[6][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][0]), 
        .b_in(b[7][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][1]), 
        .b_out(b[8][0]),
        .acc_out(d_out[7][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][1]), 
        .b_in(b[7][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][2]), 
        .b_out(b[8][1]),
        .acc_out(d_out[7][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][2]), 
        .b_in(b[7][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][3]), 
        .b_out(b[8][2]),
        .acc_out(d_out[7][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][3]), 
        .b_in(b[7][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][4]), 
        .b_out(b[8][3]),
        .acc_out(d_out[7][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][4]), 
        .b_in(b[7][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][5]), 
        .b_out(b[8][4]),
        .acc_out(d_out[7][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][5]), 
        .b_in(b[7][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][6]), 
        .b_out(b[8][5]),
        .acc_out(d_out[7][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][6]), 
        .b_in(b[7][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][7]), 
        .b_out(b[8][6]),
        .acc_out(d_out[7][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][7]), 
        .b_in(b[7][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][8]), 
        .b_out(b[8][7]),
        .acc_out(d_out[7][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][8]), 
        .b_in(b[7][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][9]), 
        .b_out(b[8][8]),
        .acc_out(d_out[7][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][9]), 
        .b_in(b[7][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][10]), 
        .b_out(b[8][9]),
        .acc_out(d_out[7][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][10]), 
        .b_in(b[7][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][11]), 
        .b_out(b[8][10]),
        .acc_out(d_out[7][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][11]), 
        .b_in(b[7][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][12]), 
        .b_out(b[8][11]),
        .acc_out(d_out[7][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][12]), 
        .b_in(b[7][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][13]), 
        .b_out(b[8][12]),
        .acc_out(d_out[7][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][13]), 
        .b_in(b[7][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][14]), 
        .b_out(b[8][13]),
        .acc_out(d_out[7][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][14]), 
        .b_in(b[7][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][15]), 
        .b_out(b[8][14]),
        .acc_out(d_out[7][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][15]), 
        .b_in(b[7][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][16]), 
        .b_out(b[8][15]),
        .acc_out(d_out[7][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][16]), 
        .b_in(b[7][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][17]), 
        .b_out(b[8][16]),
        .acc_out(d_out[7][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][17]), 
        .b_in(b[7][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][18]), 
        .b_out(b[8][17]),
        .acc_out(d_out[7][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][18]), 
        .b_in(b[7][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][19]), 
        .b_out(b[8][18]),
        .acc_out(d_out[7][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][19]), 
        .b_in(b[7][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][20]), 
        .b_out(b[8][19]),
        .acc_out(d_out[7][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][20]), 
        .b_in(b[7][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][21]), 
        .b_out(b[8][20]),
        .acc_out(d_out[7][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][21]), 
        .b_in(b[7][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][22]), 
        .b_out(b[8][21]),
        .acc_out(d_out[7][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][22]), 
        .b_in(b[7][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][23]), 
        .b_out(b[8][22]),
        .acc_out(d_out[7][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][23]), 
        .b_in(b[7][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][24]), 
        .b_out(b[8][23]),
        .acc_out(d_out[7][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][24]), 
        .b_in(b[7][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][25]), 
        .b_out(b[8][24]),
        .acc_out(d_out[7][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][25]), 
        .b_in(b[7][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][26]), 
        .b_out(b[8][25]),
        .acc_out(d_out[7][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][26]), 
        .b_in(b[7][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][27]), 
        .b_out(b[8][26]),
        .acc_out(d_out[7][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][27]), 
        .b_in(b[7][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][28]), 
        .b_out(b[8][27]),
        .acc_out(d_out[7][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][28]), 
        .b_in(b[7][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][29]), 
        .b_out(b[8][28]),
        .acc_out(d_out[7][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][29]), 
        .b_in(b[7][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][30]), 
        .b_out(b[8][29]),
        .acc_out(d_out[7][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][30]), 
        .b_in(b[7][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][31]), 
        .b_out(b[8][30]),
        .acc_out(d_out[7][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[7][31]), 
        .b_in(b[7][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[7][32]), 
        .b_out(b[8][31]),
        .acc_out(d_out[7][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][0]), 
        .b_in(b[8][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][1]), 
        .b_out(b[9][0]),
        .acc_out(d_out[8][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][1]), 
        .b_in(b[8][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][2]), 
        .b_out(b[9][1]),
        .acc_out(d_out[8][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][2]), 
        .b_in(b[8][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][3]), 
        .b_out(b[9][2]),
        .acc_out(d_out[8][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][3]), 
        .b_in(b[8][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][4]), 
        .b_out(b[9][3]),
        .acc_out(d_out[8][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][4]), 
        .b_in(b[8][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][5]), 
        .b_out(b[9][4]),
        .acc_out(d_out[8][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][5]), 
        .b_in(b[8][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][6]), 
        .b_out(b[9][5]),
        .acc_out(d_out[8][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][6]), 
        .b_in(b[8][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][7]), 
        .b_out(b[9][6]),
        .acc_out(d_out[8][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][7]), 
        .b_in(b[8][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][8]), 
        .b_out(b[9][7]),
        .acc_out(d_out[8][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][8]), 
        .b_in(b[8][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][9]), 
        .b_out(b[9][8]),
        .acc_out(d_out[8][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][9]), 
        .b_in(b[8][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][10]), 
        .b_out(b[9][9]),
        .acc_out(d_out[8][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][10]), 
        .b_in(b[8][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][11]), 
        .b_out(b[9][10]),
        .acc_out(d_out[8][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][11]), 
        .b_in(b[8][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][12]), 
        .b_out(b[9][11]),
        .acc_out(d_out[8][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][12]), 
        .b_in(b[8][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][13]), 
        .b_out(b[9][12]),
        .acc_out(d_out[8][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][13]), 
        .b_in(b[8][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][14]), 
        .b_out(b[9][13]),
        .acc_out(d_out[8][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][14]), 
        .b_in(b[8][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][15]), 
        .b_out(b[9][14]),
        .acc_out(d_out[8][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][15]), 
        .b_in(b[8][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][16]), 
        .b_out(b[9][15]),
        .acc_out(d_out[8][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][16]), 
        .b_in(b[8][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][17]), 
        .b_out(b[9][16]),
        .acc_out(d_out[8][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][17]), 
        .b_in(b[8][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][18]), 
        .b_out(b[9][17]),
        .acc_out(d_out[8][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][18]), 
        .b_in(b[8][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][19]), 
        .b_out(b[9][18]),
        .acc_out(d_out[8][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][19]), 
        .b_in(b[8][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][20]), 
        .b_out(b[9][19]),
        .acc_out(d_out[8][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][20]), 
        .b_in(b[8][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][21]), 
        .b_out(b[9][20]),
        .acc_out(d_out[8][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][21]), 
        .b_in(b[8][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][22]), 
        .b_out(b[9][21]),
        .acc_out(d_out[8][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][22]), 
        .b_in(b[8][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][23]), 
        .b_out(b[9][22]),
        .acc_out(d_out[8][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][23]), 
        .b_in(b[8][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][24]), 
        .b_out(b[9][23]),
        .acc_out(d_out[8][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][24]), 
        .b_in(b[8][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][25]), 
        .b_out(b[9][24]),
        .acc_out(d_out[8][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][25]), 
        .b_in(b[8][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][26]), 
        .b_out(b[9][25]),
        .acc_out(d_out[8][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][26]), 
        .b_in(b[8][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][27]), 
        .b_out(b[9][26]),
        .acc_out(d_out[8][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][27]), 
        .b_in(b[8][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][28]), 
        .b_out(b[9][27]),
        .acc_out(d_out[8][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][28]), 
        .b_in(b[8][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][29]), 
        .b_out(b[9][28]),
        .acc_out(d_out[8][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][29]), 
        .b_in(b[8][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][30]), 
        .b_out(b[9][29]),
        .acc_out(d_out[8][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][30]), 
        .b_in(b[8][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][31]), 
        .b_out(b[9][30]),
        .acc_out(d_out[8][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[8][31]), 
        .b_in(b[8][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[8][32]), 
        .b_out(b[9][31]),
        .acc_out(d_out[8][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][0]), 
        .b_in(b[9][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][1]), 
        .b_out(b[10][0]),
        .acc_out(d_out[9][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][1]), 
        .b_in(b[9][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][2]), 
        .b_out(b[10][1]),
        .acc_out(d_out[9][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][2]), 
        .b_in(b[9][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][3]), 
        .b_out(b[10][2]),
        .acc_out(d_out[9][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][3]), 
        .b_in(b[9][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][4]), 
        .b_out(b[10][3]),
        .acc_out(d_out[9][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][4]), 
        .b_in(b[9][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][5]), 
        .b_out(b[10][4]),
        .acc_out(d_out[9][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][5]), 
        .b_in(b[9][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][6]), 
        .b_out(b[10][5]),
        .acc_out(d_out[9][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][6]), 
        .b_in(b[9][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][7]), 
        .b_out(b[10][6]),
        .acc_out(d_out[9][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][7]), 
        .b_in(b[9][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][8]), 
        .b_out(b[10][7]),
        .acc_out(d_out[9][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][8]), 
        .b_in(b[9][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][9]), 
        .b_out(b[10][8]),
        .acc_out(d_out[9][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][9]), 
        .b_in(b[9][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][10]), 
        .b_out(b[10][9]),
        .acc_out(d_out[9][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][10]), 
        .b_in(b[9][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][11]), 
        .b_out(b[10][10]),
        .acc_out(d_out[9][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][11]), 
        .b_in(b[9][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][12]), 
        .b_out(b[10][11]),
        .acc_out(d_out[9][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][12]), 
        .b_in(b[9][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][13]), 
        .b_out(b[10][12]),
        .acc_out(d_out[9][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][13]), 
        .b_in(b[9][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][14]), 
        .b_out(b[10][13]),
        .acc_out(d_out[9][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][14]), 
        .b_in(b[9][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][15]), 
        .b_out(b[10][14]),
        .acc_out(d_out[9][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][15]), 
        .b_in(b[9][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][16]), 
        .b_out(b[10][15]),
        .acc_out(d_out[9][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][16]), 
        .b_in(b[9][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][17]), 
        .b_out(b[10][16]),
        .acc_out(d_out[9][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][17]), 
        .b_in(b[9][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][18]), 
        .b_out(b[10][17]),
        .acc_out(d_out[9][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][18]), 
        .b_in(b[9][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][19]), 
        .b_out(b[10][18]),
        .acc_out(d_out[9][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][19]), 
        .b_in(b[9][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][20]), 
        .b_out(b[10][19]),
        .acc_out(d_out[9][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][20]), 
        .b_in(b[9][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][21]), 
        .b_out(b[10][20]),
        .acc_out(d_out[9][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][21]), 
        .b_in(b[9][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][22]), 
        .b_out(b[10][21]),
        .acc_out(d_out[9][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][22]), 
        .b_in(b[9][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][23]), 
        .b_out(b[10][22]),
        .acc_out(d_out[9][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][23]), 
        .b_in(b[9][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][24]), 
        .b_out(b[10][23]),
        .acc_out(d_out[9][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][24]), 
        .b_in(b[9][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][25]), 
        .b_out(b[10][24]),
        .acc_out(d_out[9][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][25]), 
        .b_in(b[9][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][26]), 
        .b_out(b[10][25]),
        .acc_out(d_out[9][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][26]), 
        .b_in(b[9][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][27]), 
        .b_out(b[10][26]),
        .acc_out(d_out[9][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][27]), 
        .b_in(b[9][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][28]), 
        .b_out(b[10][27]),
        .acc_out(d_out[9][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][28]), 
        .b_in(b[9][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][29]), 
        .b_out(b[10][28]),
        .acc_out(d_out[9][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][29]), 
        .b_in(b[9][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][30]), 
        .b_out(b[10][29]),
        .acc_out(d_out[9][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][30]), 
        .b_in(b[9][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][31]), 
        .b_out(b[10][30]),
        .acc_out(d_out[9][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[9][31]), 
        .b_in(b[9][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[9][32]), 
        .b_out(b[10][31]),
        .acc_out(d_out[9][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][0]), 
        .b_in(b[10][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][1]), 
        .b_out(b[11][0]),
        .acc_out(d_out[10][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][1]), 
        .b_in(b[10][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][2]), 
        .b_out(b[11][1]),
        .acc_out(d_out[10][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][2]), 
        .b_in(b[10][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][3]), 
        .b_out(b[11][2]),
        .acc_out(d_out[10][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][3]), 
        .b_in(b[10][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][4]), 
        .b_out(b[11][3]),
        .acc_out(d_out[10][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][4]), 
        .b_in(b[10][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][5]), 
        .b_out(b[11][4]),
        .acc_out(d_out[10][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][5]), 
        .b_in(b[10][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][6]), 
        .b_out(b[11][5]),
        .acc_out(d_out[10][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][6]), 
        .b_in(b[10][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][7]), 
        .b_out(b[11][6]),
        .acc_out(d_out[10][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][7]), 
        .b_in(b[10][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][8]), 
        .b_out(b[11][7]),
        .acc_out(d_out[10][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][8]), 
        .b_in(b[10][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][9]), 
        .b_out(b[11][8]),
        .acc_out(d_out[10][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][9]), 
        .b_in(b[10][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][10]), 
        .b_out(b[11][9]),
        .acc_out(d_out[10][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][10]), 
        .b_in(b[10][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][11]), 
        .b_out(b[11][10]),
        .acc_out(d_out[10][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][11]), 
        .b_in(b[10][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][12]), 
        .b_out(b[11][11]),
        .acc_out(d_out[10][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][12]), 
        .b_in(b[10][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][13]), 
        .b_out(b[11][12]),
        .acc_out(d_out[10][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][13]), 
        .b_in(b[10][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][14]), 
        .b_out(b[11][13]),
        .acc_out(d_out[10][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][14]), 
        .b_in(b[10][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][15]), 
        .b_out(b[11][14]),
        .acc_out(d_out[10][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][15]), 
        .b_in(b[10][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][16]), 
        .b_out(b[11][15]),
        .acc_out(d_out[10][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][16]), 
        .b_in(b[10][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][17]), 
        .b_out(b[11][16]),
        .acc_out(d_out[10][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][17]), 
        .b_in(b[10][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][18]), 
        .b_out(b[11][17]),
        .acc_out(d_out[10][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][18]), 
        .b_in(b[10][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][19]), 
        .b_out(b[11][18]),
        .acc_out(d_out[10][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][19]), 
        .b_in(b[10][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][20]), 
        .b_out(b[11][19]),
        .acc_out(d_out[10][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][20]), 
        .b_in(b[10][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][21]), 
        .b_out(b[11][20]),
        .acc_out(d_out[10][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][21]), 
        .b_in(b[10][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][22]), 
        .b_out(b[11][21]),
        .acc_out(d_out[10][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][22]), 
        .b_in(b[10][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][23]), 
        .b_out(b[11][22]),
        .acc_out(d_out[10][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][23]), 
        .b_in(b[10][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][24]), 
        .b_out(b[11][23]),
        .acc_out(d_out[10][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][24]), 
        .b_in(b[10][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][25]), 
        .b_out(b[11][24]),
        .acc_out(d_out[10][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][25]), 
        .b_in(b[10][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][26]), 
        .b_out(b[11][25]),
        .acc_out(d_out[10][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][26]), 
        .b_in(b[10][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][27]), 
        .b_out(b[11][26]),
        .acc_out(d_out[10][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][27]), 
        .b_in(b[10][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][28]), 
        .b_out(b[11][27]),
        .acc_out(d_out[10][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][28]), 
        .b_in(b[10][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][29]), 
        .b_out(b[11][28]),
        .acc_out(d_out[10][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][29]), 
        .b_in(b[10][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][30]), 
        .b_out(b[11][29]),
        .acc_out(d_out[10][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][30]), 
        .b_in(b[10][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][31]), 
        .b_out(b[11][30]),
        .acc_out(d_out[10][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[10][31]), 
        .b_in(b[10][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[10][32]), 
        .b_out(b[11][31]),
        .acc_out(d_out[10][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][0]), 
        .b_in(b[11][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][1]), 
        .b_out(b[12][0]),
        .acc_out(d_out[11][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][1]), 
        .b_in(b[11][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][2]), 
        .b_out(b[12][1]),
        .acc_out(d_out[11][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][2]), 
        .b_in(b[11][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][3]), 
        .b_out(b[12][2]),
        .acc_out(d_out[11][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][3]), 
        .b_in(b[11][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][4]), 
        .b_out(b[12][3]),
        .acc_out(d_out[11][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][4]), 
        .b_in(b[11][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][5]), 
        .b_out(b[12][4]),
        .acc_out(d_out[11][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][5]), 
        .b_in(b[11][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][6]), 
        .b_out(b[12][5]),
        .acc_out(d_out[11][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][6]), 
        .b_in(b[11][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][7]), 
        .b_out(b[12][6]),
        .acc_out(d_out[11][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][7]), 
        .b_in(b[11][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][8]), 
        .b_out(b[12][7]),
        .acc_out(d_out[11][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][8]), 
        .b_in(b[11][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][9]), 
        .b_out(b[12][8]),
        .acc_out(d_out[11][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][9]), 
        .b_in(b[11][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][10]), 
        .b_out(b[12][9]),
        .acc_out(d_out[11][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][10]), 
        .b_in(b[11][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][11]), 
        .b_out(b[12][10]),
        .acc_out(d_out[11][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][11]), 
        .b_in(b[11][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][12]), 
        .b_out(b[12][11]),
        .acc_out(d_out[11][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][12]), 
        .b_in(b[11][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][13]), 
        .b_out(b[12][12]),
        .acc_out(d_out[11][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][13]), 
        .b_in(b[11][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][14]), 
        .b_out(b[12][13]),
        .acc_out(d_out[11][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][14]), 
        .b_in(b[11][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][15]), 
        .b_out(b[12][14]),
        .acc_out(d_out[11][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][15]), 
        .b_in(b[11][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][16]), 
        .b_out(b[12][15]),
        .acc_out(d_out[11][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][16]), 
        .b_in(b[11][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][17]), 
        .b_out(b[12][16]),
        .acc_out(d_out[11][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][17]), 
        .b_in(b[11][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][18]), 
        .b_out(b[12][17]),
        .acc_out(d_out[11][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][18]), 
        .b_in(b[11][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][19]), 
        .b_out(b[12][18]),
        .acc_out(d_out[11][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][19]), 
        .b_in(b[11][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][20]), 
        .b_out(b[12][19]),
        .acc_out(d_out[11][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][20]), 
        .b_in(b[11][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][21]), 
        .b_out(b[12][20]),
        .acc_out(d_out[11][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][21]), 
        .b_in(b[11][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][22]), 
        .b_out(b[12][21]),
        .acc_out(d_out[11][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][22]), 
        .b_in(b[11][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][23]), 
        .b_out(b[12][22]),
        .acc_out(d_out[11][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][23]), 
        .b_in(b[11][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][24]), 
        .b_out(b[12][23]),
        .acc_out(d_out[11][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][24]), 
        .b_in(b[11][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][25]), 
        .b_out(b[12][24]),
        .acc_out(d_out[11][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][25]), 
        .b_in(b[11][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][26]), 
        .b_out(b[12][25]),
        .acc_out(d_out[11][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][26]), 
        .b_in(b[11][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][27]), 
        .b_out(b[12][26]),
        .acc_out(d_out[11][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][27]), 
        .b_in(b[11][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][28]), 
        .b_out(b[12][27]),
        .acc_out(d_out[11][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][28]), 
        .b_in(b[11][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][29]), 
        .b_out(b[12][28]),
        .acc_out(d_out[11][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][29]), 
        .b_in(b[11][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][30]), 
        .b_out(b[12][29]),
        .acc_out(d_out[11][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][30]), 
        .b_in(b[11][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][31]), 
        .b_out(b[12][30]),
        .acc_out(d_out[11][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[11][31]), 
        .b_in(b[11][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[11][32]), 
        .b_out(b[12][31]),
        .acc_out(d_out[11][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][0]), 
        .b_in(b[12][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][1]), 
        .b_out(b[13][0]),
        .acc_out(d_out[12][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][1]), 
        .b_in(b[12][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][2]), 
        .b_out(b[13][1]),
        .acc_out(d_out[12][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][2]), 
        .b_in(b[12][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][3]), 
        .b_out(b[13][2]),
        .acc_out(d_out[12][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][3]), 
        .b_in(b[12][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][4]), 
        .b_out(b[13][3]),
        .acc_out(d_out[12][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][4]), 
        .b_in(b[12][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][5]), 
        .b_out(b[13][4]),
        .acc_out(d_out[12][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][5]), 
        .b_in(b[12][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][6]), 
        .b_out(b[13][5]),
        .acc_out(d_out[12][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][6]), 
        .b_in(b[12][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][7]), 
        .b_out(b[13][6]),
        .acc_out(d_out[12][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][7]), 
        .b_in(b[12][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][8]), 
        .b_out(b[13][7]),
        .acc_out(d_out[12][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][8]), 
        .b_in(b[12][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][9]), 
        .b_out(b[13][8]),
        .acc_out(d_out[12][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][9]), 
        .b_in(b[12][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][10]), 
        .b_out(b[13][9]),
        .acc_out(d_out[12][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][10]), 
        .b_in(b[12][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][11]), 
        .b_out(b[13][10]),
        .acc_out(d_out[12][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][11]), 
        .b_in(b[12][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][12]), 
        .b_out(b[13][11]),
        .acc_out(d_out[12][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][12]), 
        .b_in(b[12][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][13]), 
        .b_out(b[13][12]),
        .acc_out(d_out[12][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][13]), 
        .b_in(b[12][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][14]), 
        .b_out(b[13][13]),
        .acc_out(d_out[12][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][14]), 
        .b_in(b[12][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][15]), 
        .b_out(b[13][14]),
        .acc_out(d_out[12][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][15]), 
        .b_in(b[12][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][16]), 
        .b_out(b[13][15]),
        .acc_out(d_out[12][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][16]), 
        .b_in(b[12][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][17]), 
        .b_out(b[13][16]),
        .acc_out(d_out[12][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][17]), 
        .b_in(b[12][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][18]), 
        .b_out(b[13][17]),
        .acc_out(d_out[12][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][18]), 
        .b_in(b[12][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][19]), 
        .b_out(b[13][18]),
        .acc_out(d_out[12][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][19]), 
        .b_in(b[12][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][20]), 
        .b_out(b[13][19]),
        .acc_out(d_out[12][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][20]), 
        .b_in(b[12][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][21]), 
        .b_out(b[13][20]),
        .acc_out(d_out[12][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][21]), 
        .b_in(b[12][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][22]), 
        .b_out(b[13][21]),
        .acc_out(d_out[12][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][22]), 
        .b_in(b[12][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][23]), 
        .b_out(b[13][22]),
        .acc_out(d_out[12][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][23]), 
        .b_in(b[12][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][24]), 
        .b_out(b[13][23]),
        .acc_out(d_out[12][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][24]), 
        .b_in(b[12][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][25]), 
        .b_out(b[13][24]),
        .acc_out(d_out[12][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][25]), 
        .b_in(b[12][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][26]), 
        .b_out(b[13][25]),
        .acc_out(d_out[12][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][26]), 
        .b_in(b[12][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][27]), 
        .b_out(b[13][26]),
        .acc_out(d_out[12][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][27]), 
        .b_in(b[12][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][28]), 
        .b_out(b[13][27]),
        .acc_out(d_out[12][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][28]), 
        .b_in(b[12][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][29]), 
        .b_out(b[13][28]),
        .acc_out(d_out[12][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][29]), 
        .b_in(b[12][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][30]), 
        .b_out(b[13][29]),
        .acc_out(d_out[12][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][30]), 
        .b_in(b[12][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][31]), 
        .b_out(b[13][30]),
        .acc_out(d_out[12][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[12][31]), 
        .b_in(b[12][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[12][32]), 
        .b_out(b[13][31]),
        .acc_out(d_out[12][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][0]), 
        .b_in(b[13][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][1]), 
        .b_out(b[14][0]),
        .acc_out(d_out[13][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][1]), 
        .b_in(b[13][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][2]), 
        .b_out(b[14][1]),
        .acc_out(d_out[13][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][2]), 
        .b_in(b[13][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][3]), 
        .b_out(b[14][2]),
        .acc_out(d_out[13][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][3]), 
        .b_in(b[13][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][4]), 
        .b_out(b[14][3]),
        .acc_out(d_out[13][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][4]), 
        .b_in(b[13][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][5]), 
        .b_out(b[14][4]),
        .acc_out(d_out[13][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][5]), 
        .b_in(b[13][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][6]), 
        .b_out(b[14][5]),
        .acc_out(d_out[13][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][6]), 
        .b_in(b[13][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][7]), 
        .b_out(b[14][6]),
        .acc_out(d_out[13][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][7]), 
        .b_in(b[13][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][8]), 
        .b_out(b[14][7]),
        .acc_out(d_out[13][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][8]), 
        .b_in(b[13][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][9]), 
        .b_out(b[14][8]),
        .acc_out(d_out[13][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][9]), 
        .b_in(b[13][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][10]), 
        .b_out(b[14][9]),
        .acc_out(d_out[13][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][10]), 
        .b_in(b[13][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][11]), 
        .b_out(b[14][10]),
        .acc_out(d_out[13][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][11]), 
        .b_in(b[13][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][12]), 
        .b_out(b[14][11]),
        .acc_out(d_out[13][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][12]), 
        .b_in(b[13][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][13]), 
        .b_out(b[14][12]),
        .acc_out(d_out[13][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][13]), 
        .b_in(b[13][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][14]), 
        .b_out(b[14][13]),
        .acc_out(d_out[13][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][14]), 
        .b_in(b[13][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][15]), 
        .b_out(b[14][14]),
        .acc_out(d_out[13][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][15]), 
        .b_in(b[13][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][16]), 
        .b_out(b[14][15]),
        .acc_out(d_out[13][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][16]), 
        .b_in(b[13][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][17]), 
        .b_out(b[14][16]),
        .acc_out(d_out[13][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][17]), 
        .b_in(b[13][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][18]), 
        .b_out(b[14][17]),
        .acc_out(d_out[13][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][18]), 
        .b_in(b[13][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][19]), 
        .b_out(b[14][18]),
        .acc_out(d_out[13][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][19]), 
        .b_in(b[13][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][20]), 
        .b_out(b[14][19]),
        .acc_out(d_out[13][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][20]), 
        .b_in(b[13][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][21]), 
        .b_out(b[14][20]),
        .acc_out(d_out[13][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][21]), 
        .b_in(b[13][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][22]), 
        .b_out(b[14][21]),
        .acc_out(d_out[13][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][22]), 
        .b_in(b[13][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][23]), 
        .b_out(b[14][22]),
        .acc_out(d_out[13][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][23]), 
        .b_in(b[13][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][24]), 
        .b_out(b[14][23]),
        .acc_out(d_out[13][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][24]), 
        .b_in(b[13][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][25]), 
        .b_out(b[14][24]),
        .acc_out(d_out[13][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][25]), 
        .b_in(b[13][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][26]), 
        .b_out(b[14][25]),
        .acc_out(d_out[13][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][26]), 
        .b_in(b[13][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][27]), 
        .b_out(b[14][26]),
        .acc_out(d_out[13][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][27]), 
        .b_in(b[13][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][28]), 
        .b_out(b[14][27]),
        .acc_out(d_out[13][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][28]), 
        .b_in(b[13][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][29]), 
        .b_out(b[14][28]),
        .acc_out(d_out[13][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][29]), 
        .b_in(b[13][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][30]), 
        .b_out(b[14][29]),
        .acc_out(d_out[13][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][30]), 
        .b_in(b[13][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][31]), 
        .b_out(b[14][30]),
        .acc_out(d_out[13][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[13][31]), 
        .b_in(b[13][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[13][32]), 
        .b_out(b[14][31]),
        .acc_out(d_out[13][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][0]), 
        .b_in(b[14][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][1]), 
        .b_out(b[15][0]),
        .acc_out(d_out[14][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][1]), 
        .b_in(b[14][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][2]), 
        .b_out(b[15][1]),
        .acc_out(d_out[14][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][2]), 
        .b_in(b[14][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][3]), 
        .b_out(b[15][2]),
        .acc_out(d_out[14][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][3]), 
        .b_in(b[14][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][4]), 
        .b_out(b[15][3]),
        .acc_out(d_out[14][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][4]), 
        .b_in(b[14][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][5]), 
        .b_out(b[15][4]),
        .acc_out(d_out[14][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][5]), 
        .b_in(b[14][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][6]), 
        .b_out(b[15][5]),
        .acc_out(d_out[14][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][6]), 
        .b_in(b[14][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][7]), 
        .b_out(b[15][6]),
        .acc_out(d_out[14][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][7]), 
        .b_in(b[14][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][8]), 
        .b_out(b[15][7]),
        .acc_out(d_out[14][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][8]), 
        .b_in(b[14][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][9]), 
        .b_out(b[15][8]),
        .acc_out(d_out[14][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][9]), 
        .b_in(b[14][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][10]), 
        .b_out(b[15][9]),
        .acc_out(d_out[14][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][10]), 
        .b_in(b[14][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][11]), 
        .b_out(b[15][10]),
        .acc_out(d_out[14][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][11]), 
        .b_in(b[14][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][12]), 
        .b_out(b[15][11]),
        .acc_out(d_out[14][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][12]), 
        .b_in(b[14][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][13]), 
        .b_out(b[15][12]),
        .acc_out(d_out[14][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][13]), 
        .b_in(b[14][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][14]), 
        .b_out(b[15][13]),
        .acc_out(d_out[14][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][14]), 
        .b_in(b[14][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][15]), 
        .b_out(b[15][14]),
        .acc_out(d_out[14][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][15]), 
        .b_in(b[14][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][16]), 
        .b_out(b[15][15]),
        .acc_out(d_out[14][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][16]), 
        .b_in(b[14][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][17]), 
        .b_out(b[15][16]),
        .acc_out(d_out[14][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][17]), 
        .b_in(b[14][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][18]), 
        .b_out(b[15][17]),
        .acc_out(d_out[14][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][18]), 
        .b_in(b[14][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][19]), 
        .b_out(b[15][18]),
        .acc_out(d_out[14][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][19]), 
        .b_in(b[14][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][20]), 
        .b_out(b[15][19]),
        .acc_out(d_out[14][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][20]), 
        .b_in(b[14][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][21]), 
        .b_out(b[15][20]),
        .acc_out(d_out[14][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][21]), 
        .b_in(b[14][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][22]), 
        .b_out(b[15][21]),
        .acc_out(d_out[14][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][22]), 
        .b_in(b[14][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][23]), 
        .b_out(b[15][22]),
        .acc_out(d_out[14][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][23]), 
        .b_in(b[14][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][24]), 
        .b_out(b[15][23]),
        .acc_out(d_out[14][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][24]), 
        .b_in(b[14][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][25]), 
        .b_out(b[15][24]),
        .acc_out(d_out[14][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][25]), 
        .b_in(b[14][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][26]), 
        .b_out(b[15][25]),
        .acc_out(d_out[14][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][26]), 
        .b_in(b[14][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][27]), 
        .b_out(b[15][26]),
        .acc_out(d_out[14][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][27]), 
        .b_in(b[14][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][28]), 
        .b_out(b[15][27]),
        .acc_out(d_out[14][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][28]), 
        .b_in(b[14][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][29]), 
        .b_out(b[15][28]),
        .acc_out(d_out[14][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][29]), 
        .b_in(b[14][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][30]), 
        .b_out(b[15][29]),
        .acc_out(d_out[14][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][30]), 
        .b_in(b[14][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][31]), 
        .b_out(b[15][30]),
        .acc_out(d_out[14][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[14][31]), 
        .b_in(b[14][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[14][32]), 
        .b_out(b[15][31]),
        .acc_out(d_out[14][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][0]), 
        .b_in(b[15][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][1]), 
        .b_out(b[16][0]),
        .acc_out(d_out[15][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][1]), 
        .b_in(b[15][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][2]), 
        .b_out(b[16][1]),
        .acc_out(d_out[15][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][2]), 
        .b_in(b[15][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][3]), 
        .b_out(b[16][2]),
        .acc_out(d_out[15][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][3]), 
        .b_in(b[15][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][4]), 
        .b_out(b[16][3]),
        .acc_out(d_out[15][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][4]), 
        .b_in(b[15][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][5]), 
        .b_out(b[16][4]),
        .acc_out(d_out[15][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][5]), 
        .b_in(b[15][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][6]), 
        .b_out(b[16][5]),
        .acc_out(d_out[15][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][6]), 
        .b_in(b[15][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][7]), 
        .b_out(b[16][6]),
        .acc_out(d_out[15][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][7]), 
        .b_in(b[15][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][8]), 
        .b_out(b[16][7]),
        .acc_out(d_out[15][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][8]), 
        .b_in(b[15][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][9]), 
        .b_out(b[16][8]),
        .acc_out(d_out[15][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][9]), 
        .b_in(b[15][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][10]), 
        .b_out(b[16][9]),
        .acc_out(d_out[15][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][10]), 
        .b_in(b[15][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][11]), 
        .b_out(b[16][10]),
        .acc_out(d_out[15][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][11]), 
        .b_in(b[15][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][12]), 
        .b_out(b[16][11]),
        .acc_out(d_out[15][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][12]), 
        .b_in(b[15][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][13]), 
        .b_out(b[16][12]),
        .acc_out(d_out[15][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][13]), 
        .b_in(b[15][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][14]), 
        .b_out(b[16][13]),
        .acc_out(d_out[15][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][14]), 
        .b_in(b[15][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][15]), 
        .b_out(b[16][14]),
        .acc_out(d_out[15][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][15]), 
        .b_in(b[15][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][16]), 
        .b_out(b[16][15]),
        .acc_out(d_out[15][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][16]), 
        .b_in(b[15][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][17]), 
        .b_out(b[16][16]),
        .acc_out(d_out[15][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][17]), 
        .b_in(b[15][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][18]), 
        .b_out(b[16][17]),
        .acc_out(d_out[15][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][18]), 
        .b_in(b[15][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][19]), 
        .b_out(b[16][18]),
        .acc_out(d_out[15][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][19]), 
        .b_in(b[15][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][20]), 
        .b_out(b[16][19]),
        .acc_out(d_out[15][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][20]), 
        .b_in(b[15][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][21]), 
        .b_out(b[16][20]),
        .acc_out(d_out[15][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][21]), 
        .b_in(b[15][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][22]), 
        .b_out(b[16][21]),
        .acc_out(d_out[15][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][22]), 
        .b_in(b[15][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][23]), 
        .b_out(b[16][22]),
        .acc_out(d_out[15][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][23]), 
        .b_in(b[15][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][24]), 
        .b_out(b[16][23]),
        .acc_out(d_out[15][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][24]), 
        .b_in(b[15][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][25]), 
        .b_out(b[16][24]),
        .acc_out(d_out[15][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][25]), 
        .b_in(b[15][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][26]), 
        .b_out(b[16][25]),
        .acc_out(d_out[15][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][26]), 
        .b_in(b[15][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][27]), 
        .b_out(b[16][26]),
        .acc_out(d_out[15][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][27]), 
        .b_in(b[15][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][28]), 
        .b_out(b[16][27]),
        .acc_out(d_out[15][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][28]), 
        .b_in(b[15][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][29]), 
        .b_out(b[16][28]),
        .acc_out(d_out[15][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][29]), 
        .b_in(b[15][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][30]), 
        .b_out(b[16][29]),
        .acc_out(d_out[15][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][30]), 
        .b_in(b[15][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][31]), 
        .b_out(b[16][30]),
        .acc_out(d_out[15][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[15][31]), 
        .b_in(b[15][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[15][32]), 
        .b_out(b[16][31]),
        .acc_out(d_out[15][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][0]), 
        .b_in(b[16][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][1]), 
        .b_out(b[17][0]),
        .acc_out(d_out[16][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][1]), 
        .b_in(b[16][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][2]), 
        .b_out(b[17][1]),
        .acc_out(d_out[16][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][2]), 
        .b_in(b[16][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][3]), 
        .b_out(b[17][2]),
        .acc_out(d_out[16][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][3]), 
        .b_in(b[16][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][4]), 
        .b_out(b[17][3]),
        .acc_out(d_out[16][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][4]), 
        .b_in(b[16][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][5]), 
        .b_out(b[17][4]),
        .acc_out(d_out[16][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][5]), 
        .b_in(b[16][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][6]), 
        .b_out(b[17][5]),
        .acc_out(d_out[16][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][6]), 
        .b_in(b[16][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][7]), 
        .b_out(b[17][6]),
        .acc_out(d_out[16][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][7]), 
        .b_in(b[16][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][8]), 
        .b_out(b[17][7]),
        .acc_out(d_out[16][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][8]), 
        .b_in(b[16][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][9]), 
        .b_out(b[17][8]),
        .acc_out(d_out[16][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][9]), 
        .b_in(b[16][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][10]), 
        .b_out(b[17][9]),
        .acc_out(d_out[16][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][10]), 
        .b_in(b[16][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][11]), 
        .b_out(b[17][10]),
        .acc_out(d_out[16][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][11]), 
        .b_in(b[16][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][12]), 
        .b_out(b[17][11]),
        .acc_out(d_out[16][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][12]), 
        .b_in(b[16][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][13]), 
        .b_out(b[17][12]),
        .acc_out(d_out[16][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][13]), 
        .b_in(b[16][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][14]), 
        .b_out(b[17][13]),
        .acc_out(d_out[16][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][14]), 
        .b_in(b[16][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][15]), 
        .b_out(b[17][14]),
        .acc_out(d_out[16][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][15]), 
        .b_in(b[16][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][16]), 
        .b_out(b[17][15]),
        .acc_out(d_out[16][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][16]), 
        .b_in(b[16][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][17]), 
        .b_out(b[17][16]),
        .acc_out(d_out[16][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][17]), 
        .b_in(b[16][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][18]), 
        .b_out(b[17][17]),
        .acc_out(d_out[16][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][18]), 
        .b_in(b[16][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][19]), 
        .b_out(b[17][18]),
        .acc_out(d_out[16][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][19]), 
        .b_in(b[16][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][20]), 
        .b_out(b[17][19]),
        .acc_out(d_out[16][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][20]), 
        .b_in(b[16][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][21]), 
        .b_out(b[17][20]),
        .acc_out(d_out[16][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][21]), 
        .b_in(b[16][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][22]), 
        .b_out(b[17][21]),
        .acc_out(d_out[16][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][22]), 
        .b_in(b[16][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][23]), 
        .b_out(b[17][22]),
        .acc_out(d_out[16][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][23]), 
        .b_in(b[16][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][24]), 
        .b_out(b[17][23]),
        .acc_out(d_out[16][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][24]), 
        .b_in(b[16][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][25]), 
        .b_out(b[17][24]),
        .acc_out(d_out[16][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][25]), 
        .b_in(b[16][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][26]), 
        .b_out(b[17][25]),
        .acc_out(d_out[16][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][26]), 
        .b_in(b[16][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][27]), 
        .b_out(b[17][26]),
        .acc_out(d_out[16][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][27]), 
        .b_in(b[16][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][28]), 
        .b_out(b[17][27]),
        .acc_out(d_out[16][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][28]), 
        .b_in(b[16][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][29]), 
        .b_out(b[17][28]),
        .acc_out(d_out[16][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][29]), 
        .b_in(b[16][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][30]), 
        .b_out(b[17][29]),
        .acc_out(d_out[16][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][30]), 
        .b_in(b[16][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][31]), 
        .b_out(b[17][30]),
        .acc_out(d_out[16][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[16][31]), 
        .b_in(b[16][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[16][32]), 
        .b_out(b[17][31]),
        .acc_out(d_out[16][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][0]), 
        .b_in(b[17][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][1]), 
        .b_out(b[18][0]),
        .acc_out(d_out[17][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][1]), 
        .b_in(b[17][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][2]), 
        .b_out(b[18][1]),
        .acc_out(d_out[17][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][2]), 
        .b_in(b[17][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][3]), 
        .b_out(b[18][2]),
        .acc_out(d_out[17][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][3]), 
        .b_in(b[17][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][4]), 
        .b_out(b[18][3]),
        .acc_out(d_out[17][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][4]), 
        .b_in(b[17][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][5]), 
        .b_out(b[18][4]),
        .acc_out(d_out[17][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][5]), 
        .b_in(b[17][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][6]), 
        .b_out(b[18][5]),
        .acc_out(d_out[17][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][6]), 
        .b_in(b[17][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][7]), 
        .b_out(b[18][6]),
        .acc_out(d_out[17][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][7]), 
        .b_in(b[17][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][8]), 
        .b_out(b[18][7]),
        .acc_out(d_out[17][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][8]), 
        .b_in(b[17][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][9]), 
        .b_out(b[18][8]),
        .acc_out(d_out[17][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][9]), 
        .b_in(b[17][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][10]), 
        .b_out(b[18][9]),
        .acc_out(d_out[17][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][10]), 
        .b_in(b[17][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][11]), 
        .b_out(b[18][10]),
        .acc_out(d_out[17][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][11]), 
        .b_in(b[17][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][12]), 
        .b_out(b[18][11]),
        .acc_out(d_out[17][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][12]), 
        .b_in(b[17][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][13]), 
        .b_out(b[18][12]),
        .acc_out(d_out[17][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][13]), 
        .b_in(b[17][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][14]), 
        .b_out(b[18][13]),
        .acc_out(d_out[17][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][14]), 
        .b_in(b[17][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][15]), 
        .b_out(b[18][14]),
        .acc_out(d_out[17][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][15]), 
        .b_in(b[17][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][16]), 
        .b_out(b[18][15]),
        .acc_out(d_out[17][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][16]), 
        .b_in(b[17][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][17]), 
        .b_out(b[18][16]),
        .acc_out(d_out[17][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][17]), 
        .b_in(b[17][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][18]), 
        .b_out(b[18][17]),
        .acc_out(d_out[17][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][18]), 
        .b_in(b[17][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][19]), 
        .b_out(b[18][18]),
        .acc_out(d_out[17][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][19]), 
        .b_in(b[17][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][20]), 
        .b_out(b[18][19]),
        .acc_out(d_out[17][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][20]), 
        .b_in(b[17][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][21]), 
        .b_out(b[18][20]),
        .acc_out(d_out[17][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][21]), 
        .b_in(b[17][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][22]), 
        .b_out(b[18][21]),
        .acc_out(d_out[17][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][22]), 
        .b_in(b[17][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][23]), 
        .b_out(b[18][22]),
        .acc_out(d_out[17][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][23]), 
        .b_in(b[17][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][24]), 
        .b_out(b[18][23]),
        .acc_out(d_out[17][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][24]), 
        .b_in(b[17][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][25]), 
        .b_out(b[18][24]),
        .acc_out(d_out[17][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][25]), 
        .b_in(b[17][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][26]), 
        .b_out(b[18][25]),
        .acc_out(d_out[17][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][26]), 
        .b_in(b[17][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][27]), 
        .b_out(b[18][26]),
        .acc_out(d_out[17][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][27]), 
        .b_in(b[17][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][28]), 
        .b_out(b[18][27]),
        .acc_out(d_out[17][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][28]), 
        .b_in(b[17][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][29]), 
        .b_out(b[18][28]),
        .acc_out(d_out[17][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][29]), 
        .b_in(b[17][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][30]), 
        .b_out(b[18][29]),
        .acc_out(d_out[17][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][30]), 
        .b_in(b[17][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][31]), 
        .b_out(b[18][30]),
        .acc_out(d_out[17][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[17][31]), 
        .b_in(b[17][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[17][32]), 
        .b_out(b[18][31]),
        .acc_out(d_out[17][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][0]), 
        .b_in(b[18][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][1]), 
        .b_out(b[19][0]),
        .acc_out(d_out[18][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][1]), 
        .b_in(b[18][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][2]), 
        .b_out(b[19][1]),
        .acc_out(d_out[18][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][2]), 
        .b_in(b[18][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][3]), 
        .b_out(b[19][2]),
        .acc_out(d_out[18][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][3]), 
        .b_in(b[18][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][4]), 
        .b_out(b[19][3]),
        .acc_out(d_out[18][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][4]), 
        .b_in(b[18][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][5]), 
        .b_out(b[19][4]),
        .acc_out(d_out[18][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][5]), 
        .b_in(b[18][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][6]), 
        .b_out(b[19][5]),
        .acc_out(d_out[18][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][6]), 
        .b_in(b[18][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][7]), 
        .b_out(b[19][6]),
        .acc_out(d_out[18][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][7]), 
        .b_in(b[18][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][8]), 
        .b_out(b[19][7]),
        .acc_out(d_out[18][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][8]), 
        .b_in(b[18][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][9]), 
        .b_out(b[19][8]),
        .acc_out(d_out[18][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][9]), 
        .b_in(b[18][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][10]), 
        .b_out(b[19][9]),
        .acc_out(d_out[18][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][10]), 
        .b_in(b[18][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][11]), 
        .b_out(b[19][10]),
        .acc_out(d_out[18][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][11]), 
        .b_in(b[18][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][12]), 
        .b_out(b[19][11]),
        .acc_out(d_out[18][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][12]), 
        .b_in(b[18][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][13]), 
        .b_out(b[19][12]),
        .acc_out(d_out[18][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][13]), 
        .b_in(b[18][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][14]), 
        .b_out(b[19][13]),
        .acc_out(d_out[18][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][14]), 
        .b_in(b[18][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][15]), 
        .b_out(b[19][14]),
        .acc_out(d_out[18][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][15]), 
        .b_in(b[18][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][16]), 
        .b_out(b[19][15]),
        .acc_out(d_out[18][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][16]), 
        .b_in(b[18][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][17]), 
        .b_out(b[19][16]),
        .acc_out(d_out[18][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][17]), 
        .b_in(b[18][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][18]), 
        .b_out(b[19][17]),
        .acc_out(d_out[18][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][18]), 
        .b_in(b[18][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][19]), 
        .b_out(b[19][18]),
        .acc_out(d_out[18][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][19]), 
        .b_in(b[18][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][20]), 
        .b_out(b[19][19]),
        .acc_out(d_out[18][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][20]), 
        .b_in(b[18][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][21]), 
        .b_out(b[19][20]),
        .acc_out(d_out[18][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][21]), 
        .b_in(b[18][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][22]), 
        .b_out(b[19][21]),
        .acc_out(d_out[18][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][22]), 
        .b_in(b[18][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][23]), 
        .b_out(b[19][22]),
        .acc_out(d_out[18][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][23]), 
        .b_in(b[18][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][24]), 
        .b_out(b[19][23]),
        .acc_out(d_out[18][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][24]), 
        .b_in(b[18][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][25]), 
        .b_out(b[19][24]),
        .acc_out(d_out[18][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][25]), 
        .b_in(b[18][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][26]), 
        .b_out(b[19][25]),
        .acc_out(d_out[18][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][26]), 
        .b_in(b[18][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][27]), 
        .b_out(b[19][26]),
        .acc_out(d_out[18][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][27]), 
        .b_in(b[18][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][28]), 
        .b_out(b[19][27]),
        .acc_out(d_out[18][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][28]), 
        .b_in(b[18][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][29]), 
        .b_out(b[19][28]),
        .acc_out(d_out[18][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][29]), 
        .b_in(b[18][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][30]), 
        .b_out(b[19][29]),
        .acc_out(d_out[18][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][30]), 
        .b_in(b[18][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][31]), 
        .b_out(b[19][30]),
        .acc_out(d_out[18][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[18][31]), 
        .b_in(b[18][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[18][32]), 
        .b_out(b[19][31]),
        .acc_out(d_out[18][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][0]), 
        .b_in(b[19][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][1]), 
        .b_out(b[20][0]),
        .acc_out(d_out[19][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][1]), 
        .b_in(b[19][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][2]), 
        .b_out(b[20][1]),
        .acc_out(d_out[19][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][2]), 
        .b_in(b[19][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][3]), 
        .b_out(b[20][2]),
        .acc_out(d_out[19][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][3]), 
        .b_in(b[19][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][4]), 
        .b_out(b[20][3]),
        .acc_out(d_out[19][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][4]), 
        .b_in(b[19][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][5]), 
        .b_out(b[20][4]),
        .acc_out(d_out[19][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][5]), 
        .b_in(b[19][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][6]), 
        .b_out(b[20][5]),
        .acc_out(d_out[19][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][6]), 
        .b_in(b[19][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][7]), 
        .b_out(b[20][6]),
        .acc_out(d_out[19][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][7]), 
        .b_in(b[19][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][8]), 
        .b_out(b[20][7]),
        .acc_out(d_out[19][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][8]), 
        .b_in(b[19][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][9]), 
        .b_out(b[20][8]),
        .acc_out(d_out[19][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][9]), 
        .b_in(b[19][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][10]), 
        .b_out(b[20][9]),
        .acc_out(d_out[19][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][10]), 
        .b_in(b[19][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][11]), 
        .b_out(b[20][10]),
        .acc_out(d_out[19][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][11]), 
        .b_in(b[19][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][12]), 
        .b_out(b[20][11]),
        .acc_out(d_out[19][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][12]), 
        .b_in(b[19][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][13]), 
        .b_out(b[20][12]),
        .acc_out(d_out[19][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][13]), 
        .b_in(b[19][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][14]), 
        .b_out(b[20][13]),
        .acc_out(d_out[19][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][14]), 
        .b_in(b[19][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][15]), 
        .b_out(b[20][14]),
        .acc_out(d_out[19][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][15]), 
        .b_in(b[19][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][16]), 
        .b_out(b[20][15]),
        .acc_out(d_out[19][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][16]), 
        .b_in(b[19][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][17]), 
        .b_out(b[20][16]),
        .acc_out(d_out[19][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][17]), 
        .b_in(b[19][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][18]), 
        .b_out(b[20][17]),
        .acc_out(d_out[19][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][18]), 
        .b_in(b[19][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][19]), 
        .b_out(b[20][18]),
        .acc_out(d_out[19][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][19]), 
        .b_in(b[19][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][20]), 
        .b_out(b[20][19]),
        .acc_out(d_out[19][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][20]), 
        .b_in(b[19][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][21]), 
        .b_out(b[20][20]),
        .acc_out(d_out[19][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][21]), 
        .b_in(b[19][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][22]), 
        .b_out(b[20][21]),
        .acc_out(d_out[19][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][22]), 
        .b_in(b[19][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][23]), 
        .b_out(b[20][22]),
        .acc_out(d_out[19][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][23]), 
        .b_in(b[19][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][24]), 
        .b_out(b[20][23]),
        .acc_out(d_out[19][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][24]), 
        .b_in(b[19][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][25]), 
        .b_out(b[20][24]),
        .acc_out(d_out[19][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][25]), 
        .b_in(b[19][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][26]), 
        .b_out(b[20][25]),
        .acc_out(d_out[19][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][26]), 
        .b_in(b[19][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][27]), 
        .b_out(b[20][26]),
        .acc_out(d_out[19][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][27]), 
        .b_in(b[19][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][28]), 
        .b_out(b[20][27]),
        .acc_out(d_out[19][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][28]), 
        .b_in(b[19][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][29]), 
        .b_out(b[20][28]),
        .acc_out(d_out[19][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][29]), 
        .b_in(b[19][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][30]), 
        .b_out(b[20][29]),
        .acc_out(d_out[19][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][30]), 
        .b_in(b[19][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][31]), 
        .b_out(b[20][30]),
        .acc_out(d_out[19][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[19][31]), 
        .b_in(b[19][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[19][32]), 
        .b_out(b[20][31]),
        .acc_out(d_out[19][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][0]), 
        .b_in(b[20][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][1]), 
        .b_out(b[21][0]),
        .acc_out(d_out[20][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][1]), 
        .b_in(b[20][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][2]), 
        .b_out(b[21][1]),
        .acc_out(d_out[20][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][2]), 
        .b_in(b[20][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][3]), 
        .b_out(b[21][2]),
        .acc_out(d_out[20][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][3]), 
        .b_in(b[20][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][4]), 
        .b_out(b[21][3]),
        .acc_out(d_out[20][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][4]), 
        .b_in(b[20][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][5]), 
        .b_out(b[21][4]),
        .acc_out(d_out[20][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][5]), 
        .b_in(b[20][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][6]), 
        .b_out(b[21][5]),
        .acc_out(d_out[20][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][6]), 
        .b_in(b[20][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][7]), 
        .b_out(b[21][6]),
        .acc_out(d_out[20][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][7]), 
        .b_in(b[20][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][8]), 
        .b_out(b[21][7]),
        .acc_out(d_out[20][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][8]), 
        .b_in(b[20][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][9]), 
        .b_out(b[21][8]),
        .acc_out(d_out[20][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][9]), 
        .b_in(b[20][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][10]), 
        .b_out(b[21][9]),
        .acc_out(d_out[20][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][10]), 
        .b_in(b[20][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][11]), 
        .b_out(b[21][10]),
        .acc_out(d_out[20][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][11]), 
        .b_in(b[20][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][12]), 
        .b_out(b[21][11]),
        .acc_out(d_out[20][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][12]), 
        .b_in(b[20][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][13]), 
        .b_out(b[21][12]),
        .acc_out(d_out[20][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][13]), 
        .b_in(b[20][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][14]), 
        .b_out(b[21][13]),
        .acc_out(d_out[20][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][14]), 
        .b_in(b[20][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][15]), 
        .b_out(b[21][14]),
        .acc_out(d_out[20][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][15]), 
        .b_in(b[20][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][16]), 
        .b_out(b[21][15]),
        .acc_out(d_out[20][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][16]), 
        .b_in(b[20][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][17]), 
        .b_out(b[21][16]),
        .acc_out(d_out[20][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][17]), 
        .b_in(b[20][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][18]), 
        .b_out(b[21][17]),
        .acc_out(d_out[20][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][18]), 
        .b_in(b[20][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][19]), 
        .b_out(b[21][18]),
        .acc_out(d_out[20][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][19]), 
        .b_in(b[20][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][20]), 
        .b_out(b[21][19]),
        .acc_out(d_out[20][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][20]), 
        .b_in(b[20][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][21]), 
        .b_out(b[21][20]),
        .acc_out(d_out[20][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][21]), 
        .b_in(b[20][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][22]), 
        .b_out(b[21][21]),
        .acc_out(d_out[20][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][22]), 
        .b_in(b[20][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][23]), 
        .b_out(b[21][22]),
        .acc_out(d_out[20][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][23]), 
        .b_in(b[20][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][24]), 
        .b_out(b[21][23]),
        .acc_out(d_out[20][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][24]), 
        .b_in(b[20][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][25]), 
        .b_out(b[21][24]),
        .acc_out(d_out[20][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][25]), 
        .b_in(b[20][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][26]), 
        .b_out(b[21][25]),
        .acc_out(d_out[20][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][26]), 
        .b_in(b[20][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][27]), 
        .b_out(b[21][26]),
        .acc_out(d_out[20][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][27]), 
        .b_in(b[20][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][28]), 
        .b_out(b[21][27]),
        .acc_out(d_out[20][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][28]), 
        .b_in(b[20][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][29]), 
        .b_out(b[21][28]),
        .acc_out(d_out[20][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][29]), 
        .b_in(b[20][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][30]), 
        .b_out(b[21][29]),
        .acc_out(d_out[20][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][30]), 
        .b_in(b[20][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][31]), 
        .b_out(b[21][30]),
        .acc_out(d_out[20][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[20][31]), 
        .b_in(b[20][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[20][32]), 
        .b_out(b[21][31]),
        .acc_out(d_out[20][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][0]), 
        .b_in(b[21][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][1]), 
        .b_out(b[22][0]),
        .acc_out(d_out[21][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][1]), 
        .b_in(b[21][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][2]), 
        .b_out(b[22][1]),
        .acc_out(d_out[21][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][2]), 
        .b_in(b[21][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][3]), 
        .b_out(b[22][2]),
        .acc_out(d_out[21][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][3]), 
        .b_in(b[21][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][4]), 
        .b_out(b[22][3]),
        .acc_out(d_out[21][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][4]), 
        .b_in(b[21][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][5]), 
        .b_out(b[22][4]),
        .acc_out(d_out[21][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][5]), 
        .b_in(b[21][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][6]), 
        .b_out(b[22][5]),
        .acc_out(d_out[21][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][6]), 
        .b_in(b[21][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][7]), 
        .b_out(b[22][6]),
        .acc_out(d_out[21][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][7]), 
        .b_in(b[21][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][8]), 
        .b_out(b[22][7]),
        .acc_out(d_out[21][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][8]), 
        .b_in(b[21][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][9]), 
        .b_out(b[22][8]),
        .acc_out(d_out[21][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][9]), 
        .b_in(b[21][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][10]), 
        .b_out(b[22][9]),
        .acc_out(d_out[21][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][10]), 
        .b_in(b[21][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][11]), 
        .b_out(b[22][10]),
        .acc_out(d_out[21][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][11]), 
        .b_in(b[21][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][12]), 
        .b_out(b[22][11]),
        .acc_out(d_out[21][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][12]), 
        .b_in(b[21][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][13]), 
        .b_out(b[22][12]),
        .acc_out(d_out[21][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][13]), 
        .b_in(b[21][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][14]), 
        .b_out(b[22][13]),
        .acc_out(d_out[21][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][14]), 
        .b_in(b[21][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][15]), 
        .b_out(b[22][14]),
        .acc_out(d_out[21][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][15]), 
        .b_in(b[21][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][16]), 
        .b_out(b[22][15]),
        .acc_out(d_out[21][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][16]), 
        .b_in(b[21][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][17]), 
        .b_out(b[22][16]),
        .acc_out(d_out[21][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][17]), 
        .b_in(b[21][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][18]), 
        .b_out(b[22][17]),
        .acc_out(d_out[21][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][18]), 
        .b_in(b[21][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][19]), 
        .b_out(b[22][18]),
        .acc_out(d_out[21][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][19]), 
        .b_in(b[21][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][20]), 
        .b_out(b[22][19]),
        .acc_out(d_out[21][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][20]), 
        .b_in(b[21][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][21]), 
        .b_out(b[22][20]),
        .acc_out(d_out[21][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][21]), 
        .b_in(b[21][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][22]), 
        .b_out(b[22][21]),
        .acc_out(d_out[21][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][22]), 
        .b_in(b[21][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][23]), 
        .b_out(b[22][22]),
        .acc_out(d_out[21][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][23]), 
        .b_in(b[21][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][24]), 
        .b_out(b[22][23]),
        .acc_out(d_out[21][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][24]), 
        .b_in(b[21][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][25]), 
        .b_out(b[22][24]),
        .acc_out(d_out[21][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][25]), 
        .b_in(b[21][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][26]), 
        .b_out(b[22][25]),
        .acc_out(d_out[21][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][26]), 
        .b_in(b[21][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][27]), 
        .b_out(b[22][26]),
        .acc_out(d_out[21][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][27]), 
        .b_in(b[21][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][28]), 
        .b_out(b[22][27]),
        .acc_out(d_out[21][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][28]), 
        .b_in(b[21][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][29]), 
        .b_out(b[22][28]),
        .acc_out(d_out[21][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][29]), 
        .b_in(b[21][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][30]), 
        .b_out(b[22][29]),
        .acc_out(d_out[21][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][30]), 
        .b_in(b[21][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][31]), 
        .b_out(b[22][30]),
        .acc_out(d_out[21][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[21][31]), 
        .b_in(b[21][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[21][32]), 
        .b_out(b[22][31]),
        .acc_out(d_out[21][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][0]), 
        .b_in(b[22][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][1]), 
        .b_out(b[23][0]),
        .acc_out(d_out[22][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][1]), 
        .b_in(b[22][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][2]), 
        .b_out(b[23][1]),
        .acc_out(d_out[22][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][2]), 
        .b_in(b[22][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][3]), 
        .b_out(b[23][2]),
        .acc_out(d_out[22][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][3]), 
        .b_in(b[22][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][4]), 
        .b_out(b[23][3]),
        .acc_out(d_out[22][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][4]), 
        .b_in(b[22][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][5]), 
        .b_out(b[23][4]),
        .acc_out(d_out[22][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][5]), 
        .b_in(b[22][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][6]), 
        .b_out(b[23][5]),
        .acc_out(d_out[22][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][6]), 
        .b_in(b[22][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][7]), 
        .b_out(b[23][6]),
        .acc_out(d_out[22][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][7]), 
        .b_in(b[22][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][8]), 
        .b_out(b[23][7]),
        .acc_out(d_out[22][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][8]), 
        .b_in(b[22][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][9]), 
        .b_out(b[23][8]),
        .acc_out(d_out[22][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][9]), 
        .b_in(b[22][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][10]), 
        .b_out(b[23][9]),
        .acc_out(d_out[22][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][10]), 
        .b_in(b[22][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][11]), 
        .b_out(b[23][10]),
        .acc_out(d_out[22][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][11]), 
        .b_in(b[22][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][12]), 
        .b_out(b[23][11]),
        .acc_out(d_out[22][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][12]), 
        .b_in(b[22][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][13]), 
        .b_out(b[23][12]),
        .acc_out(d_out[22][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][13]), 
        .b_in(b[22][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][14]), 
        .b_out(b[23][13]),
        .acc_out(d_out[22][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][14]), 
        .b_in(b[22][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][15]), 
        .b_out(b[23][14]),
        .acc_out(d_out[22][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][15]), 
        .b_in(b[22][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][16]), 
        .b_out(b[23][15]),
        .acc_out(d_out[22][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][16]), 
        .b_in(b[22][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][17]), 
        .b_out(b[23][16]),
        .acc_out(d_out[22][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][17]), 
        .b_in(b[22][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][18]), 
        .b_out(b[23][17]),
        .acc_out(d_out[22][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][18]), 
        .b_in(b[22][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][19]), 
        .b_out(b[23][18]),
        .acc_out(d_out[22][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][19]), 
        .b_in(b[22][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][20]), 
        .b_out(b[23][19]),
        .acc_out(d_out[22][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][20]), 
        .b_in(b[22][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][21]), 
        .b_out(b[23][20]),
        .acc_out(d_out[22][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][21]), 
        .b_in(b[22][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][22]), 
        .b_out(b[23][21]),
        .acc_out(d_out[22][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][22]), 
        .b_in(b[22][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][23]), 
        .b_out(b[23][22]),
        .acc_out(d_out[22][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][23]), 
        .b_in(b[22][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][24]), 
        .b_out(b[23][23]),
        .acc_out(d_out[22][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][24]), 
        .b_in(b[22][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][25]), 
        .b_out(b[23][24]),
        .acc_out(d_out[22][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][25]), 
        .b_in(b[22][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][26]), 
        .b_out(b[23][25]),
        .acc_out(d_out[22][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][26]), 
        .b_in(b[22][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][27]), 
        .b_out(b[23][26]),
        .acc_out(d_out[22][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][27]), 
        .b_in(b[22][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][28]), 
        .b_out(b[23][27]),
        .acc_out(d_out[22][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][28]), 
        .b_in(b[22][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][29]), 
        .b_out(b[23][28]),
        .acc_out(d_out[22][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][29]), 
        .b_in(b[22][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][30]), 
        .b_out(b[23][29]),
        .acc_out(d_out[22][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][30]), 
        .b_in(b[22][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][31]), 
        .b_out(b[23][30]),
        .acc_out(d_out[22][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[22][31]), 
        .b_in(b[22][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[22][32]), 
        .b_out(b[23][31]),
        .acc_out(d_out[22][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][0]), 
        .b_in(b[23][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][1]), 
        .b_out(b[24][0]),
        .acc_out(d_out[23][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][1]), 
        .b_in(b[23][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][2]), 
        .b_out(b[24][1]),
        .acc_out(d_out[23][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][2]), 
        .b_in(b[23][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][3]), 
        .b_out(b[24][2]),
        .acc_out(d_out[23][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][3]), 
        .b_in(b[23][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][4]), 
        .b_out(b[24][3]),
        .acc_out(d_out[23][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][4]), 
        .b_in(b[23][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][5]), 
        .b_out(b[24][4]),
        .acc_out(d_out[23][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][5]), 
        .b_in(b[23][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][6]), 
        .b_out(b[24][5]),
        .acc_out(d_out[23][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][6]), 
        .b_in(b[23][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][7]), 
        .b_out(b[24][6]),
        .acc_out(d_out[23][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][7]), 
        .b_in(b[23][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][8]), 
        .b_out(b[24][7]),
        .acc_out(d_out[23][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][8]), 
        .b_in(b[23][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][9]), 
        .b_out(b[24][8]),
        .acc_out(d_out[23][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][9]), 
        .b_in(b[23][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][10]), 
        .b_out(b[24][9]),
        .acc_out(d_out[23][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][10]), 
        .b_in(b[23][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][11]), 
        .b_out(b[24][10]),
        .acc_out(d_out[23][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][11]), 
        .b_in(b[23][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][12]), 
        .b_out(b[24][11]),
        .acc_out(d_out[23][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][12]), 
        .b_in(b[23][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][13]), 
        .b_out(b[24][12]),
        .acc_out(d_out[23][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][13]), 
        .b_in(b[23][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][14]), 
        .b_out(b[24][13]),
        .acc_out(d_out[23][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][14]), 
        .b_in(b[23][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][15]), 
        .b_out(b[24][14]),
        .acc_out(d_out[23][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][15]), 
        .b_in(b[23][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][16]), 
        .b_out(b[24][15]),
        .acc_out(d_out[23][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][16]), 
        .b_in(b[23][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][17]), 
        .b_out(b[24][16]),
        .acc_out(d_out[23][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][17]), 
        .b_in(b[23][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][18]), 
        .b_out(b[24][17]),
        .acc_out(d_out[23][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][18]), 
        .b_in(b[23][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][19]), 
        .b_out(b[24][18]),
        .acc_out(d_out[23][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][19]), 
        .b_in(b[23][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][20]), 
        .b_out(b[24][19]),
        .acc_out(d_out[23][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][20]), 
        .b_in(b[23][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][21]), 
        .b_out(b[24][20]),
        .acc_out(d_out[23][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][21]), 
        .b_in(b[23][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][22]), 
        .b_out(b[24][21]),
        .acc_out(d_out[23][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][22]), 
        .b_in(b[23][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][23]), 
        .b_out(b[24][22]),
        .acc_out(d_out[23][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][23]), 
        .b_in(b[23][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][24]), 
        .b_out(b[24][23]),
        .acc_out(d_out[23][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][24]), 
        .b_in(b[23][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][25]), 
        .b_out(b[24][24]),
        .acc_out(d_out[23][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][25]), 
        .b_in(b[23][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][26]), 
        .b_out(b[24][25]),
        .acc_out(d_out[23][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][26]), 
        .b_in(b[23][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][27]), 
        .b_out(b[24][26]),
        .acc_out(d_out[23][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][27]), 
        .b_in(b[23][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][28]), 
        .b_out(b[24][27]),
        .acc_out(d_out[23][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][28]), 
        .b_in(b[23][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][29]), 
        .b_out(b[24][28]),
        .acc_out(d_out[23][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][29]), 
        .b_in(b[23][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][30]), 
        .b_out(b[24][29]),
        .acc_out(d_out[23][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][30]), 
        .b_in(b[23][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][31]), 
        .b_out(b[24][30]),
        .acc_out(d_out[23][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[23][31]), 
        .b_in(b[23][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[23][32]), 
        .b_out(b[24][31]),
        .acc_out(d_out[23][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][0]), 
        .b_in(b[24][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][1]), 
        .b_out(b[25][0]),
        .acc_out(d_out[24][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][1]), 
        .b_in(b[24][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][2]), 
        .b_out(b[25][1]),
        .acc_out(d_out[24][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][2]), 
        .b_in(b[24][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][3]), 
        .b_out(b[25][2]),
        .acc_out(d_out[24][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][3]), 
        .b_in(b[24][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][4]), 
        .b_out(b[25][3]),
        .acc_out(d_out[24][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][4]), 
        .b_in(b[24][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][5]), 
        .b_out(b[25][4]),
        .acc_out(d_out[24][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][5]), 
        .b_in(b[24][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][6]), 
        .b_out(b[25][5]),
        .acc_out(d_out[24][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][6]), 
        .b_in(b[24][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][7]), 
        .b_out(b[25][6]),
        .acc_out(d_out[24][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][7]), 
        .b_in(b[24][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][8]), 
        .b_out(b[25][7]),
        .acc_out(d_out[24][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][8]), 
        .b_in(b[24][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][9]), 
        .b_out(b[25][8]),
        .acc_out(d_out[24][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][9]), 
        .b_in(b[24][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][10]), 
        .b_out(b[25][9]),
        .acc_out(d_out[24][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][10]), 
        .b_in(b[24][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][11]), 
        .b_out(b[25][10]),
        .acc_out(d_out[24][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][11]), 
        .b_in(b[24][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][12]), 
        .b_out(b[25][11]),
        .acc_out(d_out[24][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][12]), 
        .b_in(b[24][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][13]), 
        .b_out(b[25][12]),
        .acc_out(d_out[24][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][13]), 
        .b_in(b[24][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][14]), 
        .b_out(b[25][13]),
        .acc_out(d_out[24][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][14]), 
        .b_in(b[24][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][15]), 
        .b_out(b[25][14]),
        .acc_out(d_out[24][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][15]), 
        .b_in(b[24][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][16]), 
        .b_out(b[25][15]),
        .acc_out(d_out[24][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][16]), 
        .b_in(b[24][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][17]), 
        .b_out(b[25][16]),
        .acc_out(d_out[24][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][17]), 
        .b_in(b[24][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][18]), 
        .b_out(b[25][17]),
        .acc_out(d_out[24][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][18]), 
        .b_in(b[24][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][19]), 
        .b_out(b[25][18]),
        .acc_out(d_out[24][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][19]), 
        .b_in(b[24][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][20]), 
        .b_out(b[25][19]),
        .acc_out(d_out[24][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][20]), 
        .b_in(b[24][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][21]), 
        .b_out(b[25][20]),
        .acc_out(d_out[24][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][21]), 
        .b_in(b[24][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][22]), 
        .b_out(b[25][21]),
        .acc_out(d_out[24][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][22]), 
        .b_in(b[24][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][23]), 
        .b_out(b[25][22]),
        .acc_out(d_out[24][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][23]), 
        .b_in(b[24][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][24]), 
        .b_out(b[25][23]),
        .acc_out(d_out[24][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][24]), 
        .b_in(b[24][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][25]), 
        .b_out(b[25][24]),
        .acc_out(d_out[24][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][25]), 
        .b_in(b[24][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][26]), 
        .b_out(b[25][25]),
        .acc_out(d_out[24][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][26]), 
        .b_in(b[24][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][27]), 
        .b_out(b[25][26]),
        .acc_out(d_out[24][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][27]), 
        .b_in(b[24][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][28]), 
        .b_out(b[25][27]),
        .acc_out(d_out[24][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][28]), 
        .b_in(b[24][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][29]), 
        .b_out(b[25][28]),
        .acc_out(d_out[24][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][29]), 
        .b_in(b[24][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][30]), 
        .b_out(b[25][29]),
        .acc_out(d_out[24][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][30]), 
        .b_in(b[24][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][31]), 
        .b_out(b[25][30]),
        .acc_out(d_out[24][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[24][31]), 
        .b_in(b[24][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[24][32]), 
        .b_out(b[25][31]),
        .acc_out(d_out[24][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][0]), 
        .b_in(b[25][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][1]), 
        .b_out(b[26][0]),
        .acc_out(d_out[25][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][1]), 
        .b_in(b[25][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][2]), 
        .b_out(b[26][1]),
        .acc_out(d_out[25][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][2]), 
        .b_in(b[25][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][3]), 
        .b_out(b[26][2]),
        .acc_out(d_out[25][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][3]), 
        .b_in(b[25][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][4]), 
        .b_out(b[26][3]),
        .acc_out(d_out[25][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][4]), 
        .b_in(b[25][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][5]), 
        .b_out(b[26][4]),
        .acc_out(d_out[25][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][5]), 
        .b_in(b[25][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][6]), 
        .b_out(b[26][5]),
        .acc_out(d_out[25][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][6]), 
        .b_in(b[25][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][7]), 
        .b_out(b[26][6]),
        .acc_out(d_out[25][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][7]), 
        .b_in(b[25][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][8]), 
        .b_out(b[26][7]),
        .acc_out(d_out[25][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][8]), 
        .b_in(b[25][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][9]), 
        .b_out(b[26][8]),
        .acc_out(d_out[25][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][9]), 
        .b_in(b[25][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][10]), 
        .b_out(b[26][9]),
        .acc_out(d_out[25][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][10]), 
        .b_in(b[25][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][11]), 
        .b_out(b[26][10]),
        .acc_out(d_out[25][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][11]), 
        .b_in(b[25][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][12]), 
        .b_out(b[26][11]),
        .acc_out(d_out[25][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][12]), 
        .b_in(b[25][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][13]), 
        .b_out(b[26][12]),
        .acc_out(d_out[25][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][13]), 
        .b_in(b[25][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][14]), 
        .b_out(b[26][13]),
        .acc_out(d_out[25][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][14]), 
        .b_in(b[25][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][15]), 
        .b_out(b[26][14]),
        .acc_out(d_out[25][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][15]), 
        .b_in(b[25][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][16]), 
        .b_out(b[26][15]),
        .acc_out(d_out[25][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][16]), 
        .b_in(b[25][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][17]), 
        .b_out(b[26][16]),
        .acc_out(d_out[25][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][17]), 
        .b_in(b[25][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][18]), 
        .b_out(b[26][17]),
        .acc_out(d_out[25][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][18]), 
        .b_in(b[25][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][19]), 
        .b_out(b[26][18]),
        .acc_out(d_out[25][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][19]), 
        .b_in(b[25][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][20]), 
        .b_out(b[26][19]),
        .acc_out(d_out[25][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][20]), 
        .b_in(b[25][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][21]), 
        .b_out(b[26][20]),
        .acc_out(d_out[25][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][21]), 
        .b_in(b[25][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][22]), 
        .b_out(b[26][21]),
        .acc_out(d_out[25][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][22]), 
        .b_in(b[25][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][23]), 
        .b_out(b[26][22]),
        .acc_out(d_out[25][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][23]), 
        .b_in(b[25][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][24]), 
        .b_out(b[26][23]),
        .acc_out(d_out[25][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][24]), 
        .b_in(b[25][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][25]), 
        .b_out(b[26][24]),
        .acc_out(d_out[25][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][25]), 
        .b_in(b[25][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][26]), 
        .b_out(b[26][25]),
        .acc_out(d_out[25][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][26]), 
        .b_in(b[25][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][27]), 
        .b_out(b[26][26]),
        .acc_out(d_out[25][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][27]), 
        .b_in(b[25][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][28]), 
        .b_out(b[26][27]),
        .acc_out(d_out[25][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][28]), 
        .b_in(b[25][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][29]), 
        .b_out(b[26][28]),
        .acc_out(d_out[25][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][29]), 
        .b_in(b[25][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][30]), 
        .b_out(b[26][29]),
        .acc_out(d_out[25][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][30]), 
        .b_in(b[25][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][31]), 
        .b_out(b[26][30]),
        .acc_out(d_out[25][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[25][31]), 
        .b_in(b[25][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[25][32]), 
        .b_out(b[26][31]),
        .acc_out(d_out[25][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][0]), 
        .b_in(b[26][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][1]), 
        .b_out(b[27][0]),
        .acc_out(d_out[26][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][1]), 
        .b_in(b[26][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][2]), 
        .b_out(b[27][1]),
        .acc_out(d_out[26][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][2]), 
        .b_in(b[26][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][3]), 
        .b_out(b[27][2]),
        .acc_out(d_out[26][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][3]), 
        .b_in(b[26][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][4]), 
        .b_out(b[27][3]),
        .acc_out(d_out[26][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][4]), 
        .b_in(b[26][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][5]), 
        .b_out(b[27][4]),
        .acc_out(d_out[26][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][5]), 
        .b_in(b[26][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][6]), 
        .b_out(b[27][5]),
        .acc_out(d_out[26][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][6]), 
        .b_in(b[26][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][7]), 
        .b_out(b[27][6]),
        .acc_out(d_out[26][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][7]), 
        .b_in(b[26][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][8]), 
        .b_out(b[27][7]),
        .acc_out(d_out[26][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][8]), 
        .b_in(b[26][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][9]), 
        .b_out(b[27][8]),
        .acc_out(d_out[26][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][9]), 
        .b_in(b[26][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][10]), 
        .b_out(b[27][9]),
        .acc_out(d_out[26][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][10]), 
        .b_in(b[26][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][11]), 
        .b_out(b[27][10]),
        .acc_out(d_out[26][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][11]), 
        .b_in(b[26][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][12]), 
        .b_out(b[27][11]),
        .acc_out(d_out[26][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][12]), 
        .b_in(b[26][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][13]), 
        .b_out(b[27][12]),
        .acc_out(d_out[26][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][13]), 
        .b_in(b[26][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][14]), 
        .b_out(b[27][13]),
        .acc_out(d_out[26][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][14]), 
        .b_in(b[26][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][15]), 
        .b_out(b[27][14]),
        .acc_out(d_out[26][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][15]), 
        .b_in(b[26][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][16]), 
        .b_out(b[27][15]),
        .acc_out(d_out[26][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][16]), 
        .b_in(b[26][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][17]), 
        .b_out(b[27][16]),
        .acc_out(d_out[26][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][17]), 
        .b_in(b[26][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][18]), 
        .b_out(b[27][17]),
        .acc_out(d_out[26][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][18]), 
        .b_in(b[26][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][19]), 
        .b_out(b[27][18]),
        .acc_out(d_out[26][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][19]), 
        .b_in(b[26][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][20]), 
        .b_out(b[27][19]),
        .acc_out(d_out[26][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][20]), 
        .b_in(b[26][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][21]), 
        .b_out(b[27][20]),
        .acc_out(d_out[26][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][21]), 
        .b_in(b[26][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][22]), 
        .b_out(b[27][21]),
        .acc_out(d_out[26][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][22]), 
        .b_in(b[26][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][23]), 
        .b_out(b[27][22]),
        .acc_out(d_out[26][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][23]), 
        .b_in(b[26][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][24]), 
        .b_out(b[27][23]),
        .acc_out(d_out[26][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][24]), 
        .b_in(b[26][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][25]), 
        .b_out(b[27][24]),
        .acc_out(d_out[26][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][25]), 
        .b_in(b[26][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][26]), 
        .b_out(b[27][25]),
        .acc_out(d_out[26][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][26]), 
        .b_in(b[26][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][27]), 
        .b_out(b[27][26]),
        .acc_out(d_out[26][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][27]), 
        .b_in(b[26][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][28]), 
        .b_out(b[27][27]),
        .acc_out(d_out[26][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][28]), 
        .b_in(b[26][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][29]), 
        .b_out(b[27][28]),
        .acc_out(d_out[26][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][29]), 
        .b_in(b[26][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][30]), 
        .b_out(b[27][29]),
        .acc_out(d_out[26][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][30]), 
        .b_in(b[26][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][31]), 
        .b_out(b[27][30]),
        .acc_out(d_out[26][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[26][31]), 
        .b_in(b[26][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[26][32]), 
        .b_out(b[27][31]),
        .acc_out(d_out[26][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][0]), 
        .b_in(b[27][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][1]), 
        .b_out(b[28][0]),
        .acc_out(d_out[27][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][1]), 
        .b_in(b[27][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][2]), 
        .b_out(b[28][1]),
        .acc_out(d_out[27][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][2]), 
        .b_in(b[27][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][3]), 
        .b_out(b[28][2]),
        .acc_out(d_out[27][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][3]), 
        .b_in(b[27][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][4]), 
        .b_out(b[28][3]),
        .acc_out(d_out[27][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][4]), 
        .b_in(b[27][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][5]), 
        .b_out(b[28][4]),
        .acc_out(d_out[27][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][5]), 
        .b_in(b[27][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][6]), 
        .b_out(b[28][5]),
        .acc_out(d_out[27][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][6]), 
        .b_in(b[27][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][7]), 
        .b_out(b[28][6]),
        .acc_out(d_out[27][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][7]), 
        .b_in(b[27][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][8]), 
        .b_out(b[28][7]),
        .acc_out(d_out[27][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][8]), 
        .b_in(b[27][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][9]), 
        .b_out(b[28][8]),
        .acc_out(d_out[27][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][9]), 
        .b_in(b[27][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][10]), 
        .b_out(b[28][9]),
        .acc_out(d_out[27][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][10]), 
        .b_in(b[27][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][11]), 
        .b_out(b[28][10]),
        .acc_out(d_out[27][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][11]), 
        .b_in(b[27][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][12]), 
        .b_out(b[28][11]),
        .acc_out(d_out[27][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][12]), 
        .b_in(b[27][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][13]), 
        .b_out(b[28][12]),
        .acc_out(d_out[27][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][13]), 
        .b_in(b[27][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][14]), 
        .b_out(b[28][13]),
        .acc_out(d_out[27][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][14]), 
        .b_in(b[27][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][15]), 
        .b_out(b[28][14]),
        .acc_out(d_out[27][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][15]), 
        .b_in(b[27][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][16]), 
        .b_out(b[28][15]),
        .acc_out(d_out[27][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][16]), 
        .b_in(b[27][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][17]), 
        .b_out(b[28][16]),
        .acc_out(d_out[27][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][17]), 
        .b_in(b[27][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][18]), 
        .b_out(b[28][17]),
        .acc_out(d_out[27][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][18]), 
        .b_in(b[27][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][19]), 
        .b_out(b[28][18]),
        .acc_out(d_out[27][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][19]), 
        .b_in(b[27][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][20]), 
        .b_out(b[28][19]),
        .acc_out(d_out[27][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][20]), 
        .b_in(b[27][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][21]), 
        .b_out(b[28][20]),
        .acc_out(d_out[27][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][21]), 
        .b_in(b[27][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][22]), 
        .b_out(b[28][21]),
        .acc_out(d_out[27][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][22]), 
        .b_in(b[27][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][23]), 
        .b_out(b[28][22]),
        .acc_out(d_out[27][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][23]), 
        .b_in(b[27][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][24]), 
        .b_out(b[28][23]),
        .acc_out(d_out[27][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][24]), 
        .b_in(b[27][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][25]), 
        .b_out(b[28][24]),
        .acc_out(d_out[27][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][25]), 
        .b_in(b[27][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][26]), 
        .b_out(b[28][25]),
        .acc_out(d_out[27][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][26]), 
        .b_in(b[27][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][27]), 
        .b_out(b[28][26]),
        .acc_out(d_out[27][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][27]), 
        .b_in(b[27][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][28]), 
        .b_out(b[28][27]),
        .acc_out(d_out[27][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][28]), 
        .b_in(b[27][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][29]), 
        .b_out(b[28][28]),
        .acc_out(d_out[27][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][29]), 
        .b_in(b[27][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][30]), 
        .b_out(b[28][29]),
        .acc_out(d_out[27][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][30]), 
        .b_in(b[27][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][31]), 
        .b_out(b[28][30]),
        .acc_out(d_out[27][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[27][31]), 
        .b_in(b[27][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[27][32]), 
        .b_out(b[28][31]),
        .acc_out(d_out[27][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][0]), 
        .b_in(b[28][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][1]), 
        .b_out(b[29][0]),
        .acc_out(d_out[28][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][1]), 
        .b_in(b[28][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][2]), 
        .b_out(b[29][1]),
        .acc_out(d_out[28][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][2]), 
        .b_in(b[28][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][3]), 
        .b_out(b[29][2]),
        .acc_out(d_out[28][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][3]), 
        .b_in(b[28][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][4]), 
        .b_out(b[29][3]),
        .acc_out(d_out[28][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][4]), 
        .b_in(b[28][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][5]), 
        .b_out(b[29][4]),
        .acc_out(d_out[28][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][5]), 
        .b_in(b[28][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][6]), 
        .b_out(b[29][5]),
        .acc_out(d_out[28][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][6]), 
        .b_in(b[28][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][7]), 
        .b_out(b[29][6]),
        .acc_out(d_out[28][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][7]), 
        .b_in(b[28][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][8]), 
        .b_out(b[29][7]),
        .acc_out(d_out[28][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][8]), 
        .b_in(b[28][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][9]), 
        .b_out(b[29][8]),
        .acc_out(d_out[28][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][9]), 
        .b_in(b[28][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][10]), 
        .b_out(b[29][9]),
        .acc_out(d_out[28][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][10]), 
        .b_in(b[28][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][11]), 
        .b_out(b[29][10]),
        .acc_out(d_out[28][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][11]), 
        .b_in(b[28][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][12]), 
        .b_out(b[29][11]),
        .acc_out(d_out[28][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][12]), 
        .b_in(b[28][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][13]), 
        .b_out(b[29][12]),
        .acc_out(d_out[28][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][13]), 
        .b_in(b[28][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][14]), 
        .b_out(b[29][13]),
        .acc_out(d_out[28][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][14]), 
        .b_in(b[28][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][15]), 
        .b_out(b[29][14]),
        .acc_out(d_out[28][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][15]), 
        .b_in(b[28][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][16]), 
        .b_out(b[29][15]),
        .acc_out(d_out[28][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][16]), 
        .b_in(b[28][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][17]), 
        .b_out(b[29][16]),
        .acc_out(d_out[28][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][17]), 
        .b_in(b[28][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][18]), 
        .b_out(b[29][17]),
        .acc_out(d_out[28][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][18]), 
        .b_in(b[28][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][19]), 
        .b_out(b[29][18]),
        .acc_out(d_out[28][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][19]), 
        .b_in(b[28][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][20]), 
        .b_out(b[29][19]),
        .acc_out(d_out[28][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][20]), 
        .b_in(b[28][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][21]), 
        .b_out(b[29][20]),
        .acc_out(d_out[28][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][21]), 
        .b_in(b[28][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][22]), 
        .b_out(b[29][21]),
        .acc_out(d_out[28][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][22]), 
        .b_in(b[28][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][23]), 
        .b_out(b[29][22]),
        .acc_out(d_out[28][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][23]), 
        .b_in(b[28][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][24]), 
        .b_out(b[29][23]),
        .acc_out(d_out[28][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][24]), 
        .b_in(b[28][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][25]), 
        .b_out(b[29][24]),
        .acc_out(d_out[28][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][25]), 
        .b_in(b[28][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][26]), 
        .b_out(b[29][25]),
        .acc_out(d_out[28][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][26]), 
        .b_in(b[28][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][27]), 
        .b_out(b[29][26]),
        .acc_out(d_out[28][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][27]), 
        .b_in(b[28][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][28]), 
        .b_out(b[29][27]),
        .acc_out(d_out[28][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][28]), 
        .b_in(b[28][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][29]), 
        .b_out(b[29][28]),
        .acc_out(d_out[28][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][29]), 
        .b_in(b[28][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][30]), 
        .b_out(b[29][29]),
        .acc_out(d_out[28][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][30]), 
        .b_in(b[28][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][31]), 
        .b_out(b[29][30]),
        .acc_out(d_out[28][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[28][31]), 
        .b_in(b[28][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[28][32]), 
        .b_out(b[29][31]),
        .acc_out(d_out[28][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][0]), 
        .b_in(b[29][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][1]), 
        .b_out(b[30][0]),
        .acc_out(d_out[29][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][1]), 
        .b_in(b[29][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][2]), 
        .b_out(b[30][1]),
        .acc_out(d_out[29][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][2]), 
        .b_in(b[29][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][3]), 
        .b_out(b[30][2]),
        .acc_out(d_out[29][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][3]), 
        .b_in(b[29][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][4]), 
        .b_out(b[30][3]),
        .acc_out(d_out[29][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][4]), 
        .b_in(b[29][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][5]), 
        .b_out(b[30][4]),
        .acc_out(d_out[29][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][5]), 
        .b_in(b[29][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][6]), 
        .b_out(b[30][5]),
        .acc_out(d_out[29][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][6]), 
        .b_in(b[29][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][7]), 
        .b_out(b[30][6]),
        .acc_out(d_out[29][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][7]), 
        .b_in(b[29][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][8]), 
        .b_out(b[30][7]),
        .acc_out(d_out[29][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][8]), 
        .b_in(b[29][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][9]), 
        .b_out(b[30][8]),
        .acc_out(d_out[29][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][9]), 
        .b_in(b[29][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][10]), 
        .b_out(b[30][9]),
        .acc_out(d_out[29][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][10]), 
        .b_in(b[29][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][11]), 
        .b_out(b[30][10]),
        .acc_out(d_out[29][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][11]), 
        .b_in(b[29][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][12]), 
        .b_out(b[30][11]),
        .acc_out(d_out[29][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][12]), 
        .b_in(b[29][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][13]), 
        .b_out(b[30][12]),
        .acc_out(d_out[29][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][13]), 
        .b_in(b[29][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][14]), 
        .b_out(b[30][13]),
        .acc_out(d_out[29][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][14]), 
        .b_in(b[29][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][15]), 
        .b_out(b[30][14]),
        .acc_out(d_out[29][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][15]), 
        .b_in(b[29][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][16]), 
        .b_out(b[30][15]),
        .acc_out(d_out[29][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][16]), 
        .b_in(b[29][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][17]), 
        .b_out(b[30][16]),
        .acc_out(d_out[29][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][17]), 
        .b_in(b[29][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][18]), 
        .b_out(b[30][17]),
        .acc_out(d_out[29][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][18]), 
        .b_in(b[29][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][19]), 
        .b_out(b[30][18]),
        .acc_out(d_out[29][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][19]), 
        .b_in(b[29][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][20]), 
        .b_out(b[30][19]),
        .acc_out(d_out[29][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][20]), 
        .b_in(b[29][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][21]), 
        .b_out(b[30][20]),
        .acc_out(d_out[29][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][21]), 
        .b_in(b[29][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][22]), 
        .b_out(b[30][21]),
        .acc_out(d_out[29][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][22]), 
        .b_in(b[29][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][23]), 
        .b_out(b[30][22]),
        .acc_out(d_out[29][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][23]), 
        .b_in(b[29][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][24]), 
        .b_out(b[30][23]),
        .acc_out(d_out[29][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][24]), 
        .b_in(b[29][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][25]), 
        .b_out(b[30][24]),
        .acc_out(d_out[29][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][25]), 
        .b_in(b[29][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][26]), 
        .b_out(b[30][25]),
        .acc_out(d_out[29][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][26]), 
        .b_in(b[29][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][27]), 
        .b_out(b[30][26]),
        .acc_out(d_out[29][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][27]), 
        .b_in(b[29][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][28]), 
        .b_out(b[30][27]),
        .acc_out(d_out[29][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][28]), 
        .b_in(b[29][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][29]), 
        .b_out(b[30][28]),
        .acc_out(d_out[29][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][29]), 
        .b_in(b[29][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][30]), 
        .b_out(b[30][29]),
        .acc_out(d_out[29][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][30]), 
        .b_in(b[29][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][31]), 
        .b_out(b[30][30]),
        .acc_out(d_out[29][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[29][31]), 
        .b_in(b[29][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[29][32]), 
        .b_out(b[30][31]),
        .acc_out(d_out[29][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][0]), 
        .b_in(b[30][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][1]), 
        .b_out(b[31][0]),
        .acc_out(d_out[30][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][1]), 
        .b_in(b[30][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][2]), 
        .b_out(b[31][1]),
        .acc_out(d_out[30][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][2]), 
        .b_in(b[30][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][3]), 
        .b_out(b[31][2]),
        .acc_out(d_out[30][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][3]), 
        .b_in(b[30][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][4]), 
        .b_out(b[31][3]),
        .acc_out(d_out[30][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][4]), 
        .b_in(b[30][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][5]), 
        .b_out(b[31][4]),
        .acc_out(d_out[30][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][5]), 
        .b_in(b[30][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][6]), 
        .b_out(b[31][5]),
        .acc_out(d_out[30][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][6]), 
        .b_in(b[30][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][7]), 
        .b_out(b[31][6]),
        .acc_out(d_out[30][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][7]), 
        .b_in(b[30][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][8]), 
        .b_out(b[31][7]),
        .acc_out(d_out[30][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][8]), 
        .b_in(b[30][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][9]), 
        .b_out(b[31][8]),
        .acc_out(d_out[30][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][9]), 
        .b_in(b[30][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][10]), 
        .b_out(b[31][9]),
        .acc_out(d_out[30][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][10]), 
        .b_in(b[30][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][11]), 
        .b_out(b[31][10]),
        .acc_out(d_out[30][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][11]), 
        .b_in(b[30][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][12]), 
        .b_out(b[31][11]),
        .acc_out(d_out[30][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][12]), 
        .b_in(b[30][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][13]), 
        .b_out(b[31][12]),
        .acc_out(d_out[30][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][13]), 
        .b_in(b[30][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][14]), 
        .b_out(b[31][13]),
        .acc_out(d_out[30][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][14]), 
        .b_in(b[30][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][15]), 
        .b_out(b[31][14]),
        .acc_out(d_out[30][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][15]), 
        .b_in(b[30][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][16]), 
        .b_out(b[31][15]),
        .acc_out(d_out[30][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][16]), 
        .b_in(b[30][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][17]), 
        .b_out(b[31][16]),
        .acc_out(d_out[30][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][17]), 
        .b_in(b[30][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][18]), 
        .b_out(b[31][17]),
        .acc_out(d_out[30][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][18]), 
        .b_in(b[30][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][19]), 
        .b_out(b[31][18]),
        .acc_out(d_out[30][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][19]), 
        .b_in(b[30][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][20]), 
        .b_out(b[31][19]),
        .acc_out(d_out[30][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][20]), 
        .b_in(b[30][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][21]), 
        .b_out(b[31][20]),
        .acc_out(d_out[30][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][21]), 
        .b_in(b[30][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][22]), 
        .b_out(b[31][21]),
        .acc_out(d_out[30][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][22]), 
        .b_in(b[30][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][23]), 
        .b_out(b[31][22]),
        .acc_out(d_out[30][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][23]), 
        .b_in(b[30][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][24]), 
        .b_out(b[31][23]),
        .acc_out(d_out[30][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][24]), 
        .b_in(b[30][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][25]), 
        .b_out(b[31][24]),
        .acc_out(d_out[30][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][25]), 
        .b_in(b[30][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][26]), 
        .b_out(b[31][25]),
        .acc_out(d_out[30][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][26]), 
        .b_in(b[30][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][27]), 
        .b_out(b[31][26]),
        .acc_out(d_out[30][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][27]), 
        .b_in(b[30][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][28]), 
        .b_out(b[31][27]),
        .acc_out(d_out[30][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][28]), 
        .b_in(b[30][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][29]), 
        .b_out(b[31][28]),
        .acc_out(d_out[30][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][29]), 
        .b_in(b[30][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][30]), 
        .b_out(b[31][29]),
        .acc_out(d_out[30][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][30]), 
        .b_in(b[30][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][31]), 
        .b_out(b[31][30]),
        .acc_out(d_out[30][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[30][31]), 
        .b_in(b[30][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[30][32]), 
        .b_out(b[31][31]),
        .acc_out(d_out[30][31])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][0]), 
        .b_in(b[31][0]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][1]), 
        .b_out(b[32][0]),
        .acc_out(d_out[31][0])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][1]), 
        .b_in(b[31][1]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][2]), 
        .b_out(b[32][1]),
        .acc_out(d_out[31][1])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][2]), 
        .b_in(b[31][2]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][3]), 
        .b_out(b[32][2]),
        .acc_out(d_out[31][2])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][3]), 
        .b_in(b[31][3]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][4]), 
        .b_out(b[32][3]),
        .acc_out(d_out[31][3])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][4]), 
        .b_in(b[31][4]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][5]), 
        .b_out(b[32][4]),
        .acc_out(d_out[31][4])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][5]), 
        .b_in(b[31][5]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][6]), 
        .b_out(b[32][5]),
        .acc_out(d_out[31][5])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][6]), 
        .b_in(b[31][6]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][7]), 
        .b_out(b[32][6]),
        .acc_out(d_out[31][6])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][7]), 
        .b_in(b[31][7]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][8]), 
        .b_out(b[32][7]),
        .acc_out(d_out[31][7])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][8]), 
        .b_in(b[31][8]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][9]), 
        .b_out(b[32][8]),
        .acc_out(d_out[31][8])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][9]), 
        .b_in(b[31][9]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][10]), 
        .b_out(b[32][9]),
        .acc_out(d_out[31][9])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][10]), 
        .b_in(b[31][10]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][11]), 
        .b_out(b[32][10]),
        .acc_out(d_out[31][10])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][11]), 
        .b_in(b[31][11]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][12]), 
        .b_out(b[32][11]),
        .acc_out(d_out[31][11])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][12]), 
        .b_in(b[31][12]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][13]), 
        .b_out(b[32][12]),
        .acc_out(d_out[31][12])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][13]), 
        .b_in(b[31][13]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][14]), 
        .b_out(b[32][13]),
        .acc_out(d_out[31][13])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][14]), 
        .b_in(b[31][14]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][15]), 
        .b_out(b[32][14]),
        .acc_out(d_out[31][14])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][15]), 
        .b_in(b[31][15]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][16]), 
        .b_out(b[32][15]),
        .acc_out(d_out[31][15])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][16]), 
        .b_in(b[31][16]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][17]), 
        .b_out(b[32][16]),
        .acc_out(d_out[31][16])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][17]), 
        .b_in(b[31][17]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][18]), 
        .b_out(b[32][17]),
        .acc_out(d_out[31][17])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][18]), 
        .b_in(b[31][18]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][19]), 
        .b_out(b[32][18]),
        .acc_out(d_out[31][18])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][19]), 
        .b_in(b[31][19]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][20]), 
        .b_out(b[32][19]),
        .acc_out(d_out[31][19])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][20]), 
        .b_in(b[31][20]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][21]), 
        .b_out(b[32][20]),
        .acc_out(d_out[31][20])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][21]), 
        .b_in(b[31][21]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][22]), 
        .b_out(b[32][21]),
        .acc_out(d_out[31][21])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][22]), 
        .b_in(b[31][22]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][23]), 
        .b_out(b[32][22]),
        .acc_out(d_out[31][22])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][23]), 
        .b_in(b[31][23]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][24]), 
        .b_out(b[32][23]),
        .acc_out(d_out[31][23])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][24]), 
        .b_in(b[31][24]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][25]), 
        .b_out(b[32][24]),
        .acc_out(d_out[31][24])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][25]), 
        .b_in(b[31][25]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][26]), 
        .b_out(b[32][25]),
        .acc_out(d_out[31][25])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][26]), 
        .b_in(b[31][26]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][27]), 
        .b_out(b[32][26]),
        .acc_out(d_out[31][26])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][27]), 
        .b_in(b[31][27]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][28]), 
        .b_out(b[32][27]),
        .acc_out(d_out[31][27])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][28]), 
        .b_in(b[31][28]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][29]), 
        .b_out(b[32][28]),
        .acc_out(d_out[31][28])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][29]), 
        .b_in(b[31][29]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][30]), 
        .b_out(b[32][29]),
        .acc_out(d_out[31][29])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][30]), 
        .b_in(b[31][30]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][31]), 
        .b_out(b[32][30]),
        .acc_out(d_out[31][30])
        );

    ast_mac_v element ( 
        .clk(clk), 
        .reset(reset), 
        .a_in(a[31][31]), 
        .b_in(b[31][31]), 
        .mult_en(mult_en), 
        .acc_en(acc_en), 
        .load_en(load_en), 
        .a_out(a[31][32]), 
        .b_out(b[32][31]),
        .acc_out(d_out[31][31])
        );
endmodule
